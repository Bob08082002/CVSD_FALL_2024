package dat_0;
integer pat_num = 0;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h03776113851a475bdd6618bbbaa350d46ca40c8b12daea4f517ec7582efce78d75799334cdd14bf7705f79fed6483855d684ae04cc42e5a661558ba4938e812013728b836b75b41f57a4c882df63aec6d7d55bc0fa1b7f67d24439fbbb63edb8;
reg [511:0] golden_data = 512'h551b8a12d39ef45b066a4948a94f1ddad0942cb0c2e532d8556789ebc8dc64182627b3939256128eff6abe1c2736d702e7ff7fe499fc221d3ee2f5ec074371fe;
endpackage
package dat_1;
integer pat_num = 1;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h30baf25c570c3c70400b8f88e37ec81cd95e960bd0ffffc94bced6cdce3dfa3154e26cf2abc372e8505634d786db92d7ab5727e4048fff2519d6087634ed6d761eb9fa1ba71cadbc99ade8aa029a1f632f20442c52592e7a6c94ad3dd212768a;
reg [511:0] golden_data = 512'h5c3eff352afe1f1a9f1695fe02db6e3c76672a50ddce81c8fbaf3538eb51838e0d0ecdb5eb66d572b86f02522faac09958e705ac4fae3a5dab4ee6efab0554c0;
endpackage
package dat_2;
integer pat_num = 2;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h30998afabebf77b58b78727eef92071bbd52821a3c1bf5163c3002b7ab25ba61764163870e3872612ea8798e34c76bbf626597c72db644b6faa44b211a33a40776a07f270df7630b73a202e97828bc2780743fa30f1912529ae858cd90693134;
reg [511:0] golden_data = 512'h0be5a67cfad502fa1b25ddf2d6915b48672ad69452de0c61122d87ef941d5ba41c7eee54c460121614c396ba2d5cc5858a14416d45f5ed2d8eb9e6d58b310cac;
endpackage
package dat_3;
integer pat_num = 3;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2dc5a50d50545d291803d51753a9938c637b962bfff5076ecb4cfc43b523a1ec029a187043e22450b5f36ddfcf0a02cbb0ec26374e1e5bb61cddd32d3f326bef757b7095497020f5877048fb7fae78b193efe9cb9e82abfe02b0dfec38d32661;
reg [511:0] golden_data = 512'h6bb57eb5f16f3d6ec144938773484b079f741031b2814f26db0dea80e5bdb0502f153d28678c55689e5bfab60f14170657e3543838f6be2005cd4f1aa5ec43d4;
endpackage
package dat_4;
integer pat_num = 4;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h12942e3413f8c35864cdc9b0ec97853da5706e07d6ff7a970d6a9f919fd4dc43594c40a07c63db1e7cd870d13bab90f42ffb7813efa9b6391c79dd721d813c777086660eb384c2c8b3138a5190bbff75118d90b644d75a286d68f631dbf5a529;
reg [511:0] golden_data = 512'h44fb6259cce0f5536b353fbb1c0ef04bee7a1af248b0d4f8768b356320be1e56456c25b5f7dc5e3dca0a2dba10e4ea7f5176299ce1416796e25f1610fcb10b54;
endpackage
package dat_5;
integer pat_num = 5;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7d8b1e205f06cc13d95550364986415a87d7ece3bdd167f4908671a87fa8b711657a842790b93ea1ebd500b28d2b974bbd44e98aa0ebf558f7060d6f4ba202e41e553d4deb4310c6c7968eae5f640c83a51ed7e5be1154445eb74b3775d66dc8;
reg [511:0] golden_data = 512'h18d97e79448d559e8ee18e2b22660925c395cf71c0854437eea8f92ba1ed92e600da589d312de39cf9225789e77bbc121d0f73ebc05c1af216e818c2ec94f714;
endpackage
package dat_6;
integer pat_num = 6;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h74c3f5ff5835737c7eec648dbe20bbadbb74e4f906971196b0c6093076999f3667bbe2e83f81fe4dc2b9e859603ad2cb34eedf699e6986a59e9ed082fead67c44c783b20a28696e09b8c4b38ef290376a2fde82ca317508c7a83740b29bdd324;
reg [511:0] golden_data = 512'h62de2060f99fb24388981f93157e8d7249ffd6c133840cbd58826759af843fc26a5c9eddbc4dc39633508d0f6280a5f07b1091fbc7612013da07697dda36f198;
endpackage
package dat_7;
integer pat_num = 7;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5554f5469b35235836c99571f6d2f8802d956be8f8bb3c9f2b71dd2c24a9a6d13c18f9d11bd9d6b77ed18d68b452dc99e9c8766a90ba88aeca0d864e25170fef77f058e19385550e4c46ea6f46bbaf5ad9df8539c207fd834a67fa77a1eb830d;
reg [511:0] golden_data = 512'h392ffc3ef0d747e18be979c08bbc53467410e884e3072a9b4c7f05a2dad25fd02e6d7230890e6a66af6510438de6fec23922284933ea0e724e0a7e6135ce7de6;
endpackage
package dat_8;
integer pat_num = 8;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6fc3cd5ebcb19983b367129e145a8b3fa3472a368835aa395ae394ffd5ceb91135149150ec76ae3735a34b2c0a5ea4d27a6a6c5706476d48c4d217fe86445f981c8fd5e1c8745d9de133a3438d63174fa8ce697484c4bc1cfe489ea4ecd06e6e;
reg [511:0] golden_data = 512'h7fad666799e859620c59255e0fced3de2af3a3f0ba0f0b421d7bd8b9cc7ef32a5e1b6ee0f4c52a603ddb8a78e5a13fe1ea58ae1ff9a9932cca62d3d726d4c6bc;
endpackage
package dat_9;
integer pat_num = 9;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4ec6b3c71a6d5ee1599175830563512cdb01c2962517c8a6650ad069b8b2656f5b69b320c9c9694a5591d9c9ecc8bb40730c54880a6e26d3ec8be0ecbf040ac7666cc2ad2414da81898e133160666cd7bfc533ecb61640c44775b84a364c2a19;
reg [511:0] golden_data = 512'h2a9de38ca59a29ef95561564852b3415bec1b863211577d8511dcd77a151d602505aad365e48f51f12ef81b85cc75e8f0dc3edcea9c6315b4fa1044509e411d2;
endpackage
package dat_10;
integer pat_num = 10;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h38500f067fc004ceefb280678d0a6bc4efea682749d5b549946b35c5d0b7544c04ada0f4e80b84472a05ff1eb339af28508e670c6e30a7729aa7e3200b8df63e35dad8bcadc3e203c18effd3ec41dc44f2f5924cbc3ebf6eee4a44284afdc8de;
reg [511:0] golden_data = 512'h3e95fa9334eed830883524b37c919c797facb0e724faca43c62c7954b350be6e6bdffafe194846f5e9628c28270e868cada0ddbaec339f6e2fb0543bd59a4826;
endpackage
package dat_11;
integer pat_num = 11;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1181074f84ce6c622f995b4b18617bf15090a9f3c24b431b6e097418a3fa885f2f2629df754c04358e1b1923e3d21b55246c87b05f2bb4dbc779dddb54520fe23822203103c29d46ad4d8e68e1e3caf299bd344b99835513e532b5b0bacfdf30;
reg [511:0] golden_data = 512'h3ca9e6ae7238c99d08b7dd835e8bdf9a8fd643b475e71f8dcedd0db12902b6dc132ab6361575edafddb19f1d2ab1df0b9b9a262df1cfa322b92de5cf8652d5e4;
endpackage
package dat_12;
integer pat_num = 12;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h30f385e6badb85b7b7a57a7a3d29c0a04695d2cd204a6a708d350e28aea0dd0e65b2bcbb0a2740dc2a24c726506f176ed297545dc4cb31a0802715c2dcf9aaba510f90535161f5c09bb8e73735c2a4839dd9041a220fea02b336bc4cf5c307b8;
reg [511:0] golden_data = 512'h2b78ccd23353d84b5422fab773df88fcc7f89370b1f639716b9e41325ed8ca506a1ffa6f0e27844d0094346d9ac2d35583e69c0d86a4ffc65da1bea936d0f646;
endpackage
package dat_13;
integer pat_num = 13;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h16120a5d0af4ec8667f60856495ae7eacde0e1fd166e371cec18e642d74a0ac72433757e100ed6a296a0b802c0752ec6dfe6613665ed63c6eb1fcccce0871a5103a0550e9363c14a61ba1082c06f3acd2bb6df398e9765af036e68e58705bda2;
reg [511:0] golden_data = 512'h5ae8ae5effd1a74c63141e4fb9004e53b83b3927db29f760b0b086a3c0ff8b8418b95a4f1704963f6f2d71653bff23bb491c47f7a95201766431413360ccb22e;
endpackage
package dat_14;
integer pat_num = 14;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5f0e896c31bbec87b10538a9a96d8b3cecf892d92652ca92596d560ecb8cc0e21c69b8f8defbb7bb43449fb64a886beaaae389e3aad9bded4a816bad85f875731d2c9552c6112b7adf9217924fea8a994f65f36a0d3fdcb6abfa365cc2e5f2bf;
reg [511:0] golden_data = 512'h35cb2a156377849183b93094971ad5aeb39f60eee8512b3896623c726cb0e6983a96c74c18b520fdb9b9b750469bd1b90e48eced105b5e2b652ebe90752eccee;
endpackage
package dat_15;
integer pat_num = 15;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h444c180115e040f5d96484ab4374c68bbff6f18dd0b1b107d3d3d8c5be00097f48febb4e3df3002b0ed2f8d019fa767184d6f755966bd71e5d3ba4c3d3fadfcf77a5266455cd3ad626e3bfb7afb38946e509057e8ea01677430ad6365557485f;
reg [511:0] golden_data = 512'h4b7053aa2769e502f77759de6e66b54a10b2eda8a8c8271b7ad5bc0e1721a6ec367005bb78553e8aa9faf4b0f3b5997d126de789ceda9b83c7db613771b22124;
endpackage
package dat_16;
integer pat_num = 16;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h016925c3af865a9ddf3dc41be1f036a6df46b89a3f3b9f49258baecb3694752f6813d75ab20dc7a160b7855e8c31b59a2cfc416e1554fc29dc4daf22add4dff518f9189e5a026bf83695ea4de0f5b2650e7da539167499770ed71c26bb0abc22;
reg [511:0] golden_data = 512'h4de0ccf769d6dc7bc8e55b18e033b6e546c96e6134e986196daad5e325d2da6a0f6966ccc651c7d6ea03a6f457127d95b6a08a28a001801afdb806e231015a34;
endpackage
package dat_17;
integer pat_num = 17;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6ef427d7e578f92e3ba569e8ebdea208b9be8d6fdb83d3a0706d3210f3c442f143f5f48f439ad7d1f6729bccaa3b5ba9624ced0bad29cfac3311fd1e11a4b6f36fb6c397931caf21fbe6466dde46ebfa122e5c6cf8411a1b3f576b1f44d6b71e;
reg [511:0] golden_data = 512'h79854288ea12482cbf7c903d6f41f744542bc7cfb8ad3acfe91756d5b526ca82319d0a040dbb6def30ba9f7c30efc32c82d97e5444b006ca829209bb4ba82ade;
endpackage
package dat_18;
integer pat_num = 18;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4f359f78e119c1e7ef9794632744f60aa27689c36aeef8dad757edb48e5f2e3517452dd79b35f5aeeafce100df93ac50583da672be3a44d5c89ffd0f6ce64c856d3505bec9cf0a2aa078675d7f84c2f508fbebdded0a97a8ac4fe2c0715b8bee;
reg [511:0] golden_data = 512'h2e442adb7ee2947f1e4e82e76618aecd804e05b69244b50c64a92968fcd256e01cb373cdcfecd0be6ee48b9e4bbed308fdb8747c750d4cf5ab08b5192ce2dca8;
endpackage
package dat_19;
integer pat_num = 19;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h64ed655b4068ab910d83f867ef7cdef7fa0976da4e985371ceb1fa0b856720a63cde75635cdefa088f6ddcc65c428c6a2d6f14c486f185b289412de70095ea5c6ef085cb050c957c1838fa8864830bbb38c6e7fe155492928a8a44ad35f8f37f;
reg [511:0] golden_data = 512'h791e1916573287d3e5ffb3bf9cb3b4ce0592caec7aff0e4628b75e2e399f40fe718eb05ff162071f38f5d7ed59dfe12744ce94d4b8ce38f03dd5b25a4bad3620;
endpackage
package dat_20;
integer pat_num = 20;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h38bd2f516707cc1ba61d68a365ad0aa0cdb3f03c414ed31d889ae4558eb5fd09457731a45f8c23b0f280982e6fb142f77334b9d0aa853ae810a8410800ff3a6f6d8faeb3d6ef903b607087caca1ba53fb04b87d7e595409e433be039a42f53d6;
reg [511:0] golden_data = 512'h3900e7b210cd2246ca4a6ec72813dd0ce529ca25fc6e27e81473f7e1cbd1576243ac16c9e9821f3e999f7f7ee95dafb20c68bd837065230e283534e76a4d13da;
endpackage
package dat_21;
integer pat_num = 21;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h47d0f501b70b1e742851c1c2ec4222c5d16f3f630fb9f6c7f514aa0198bf469a1d52df3b35e7665af52f70e415bf4deb3fa876da5b9ec0282d5c0734cebf7b77721e641c54786966be2a8fa2da5c372364233b18e4dba21c495d849a8aba6949;
reg [511:0] golden_data = 512'h6b2d812e8f8e7b5740728dd35013de65e51e6ec624bb969d568c89e226a930502010715527044875a9c764318f8d0a1e0d16d352591514b47f39409ca202303a;
endpackage
package dat_22;
integer pat_num = 22;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7780d7f0a8c58eed5d483016a847b7bb7dc4fffe00b4824e0b835062fb211cf566effaccf6170e98f9335cff5ee3ad2e3430eebaa731d24a4065786d659a28b54b843ee2a0d313324a991e9a3b8d31a27589b57a701cc13ea1517a66377a5974;
reg [511:0] golden_data = 512'h683aa1a28fdd2c6bdc1f923f31d614b1befc883a00942b6064d5471587159dbc4691f24b2cd988fecf1cc001196583a8a2489e74ab450fe333ff84175600d5f6;
endpackage
package dat_23;
integer pat_num = 23;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h009aed3af4356ab56385bdace3ac0edc8c9593219e35daf7e0d9069cb14f0c7734a012f907611f22324d2a898d425cd763bdeb574475713aa3501568b85f741451bf9768bd0fa746bd09fab230388612181bf315b3b56c9f25e7cdc64a9290d1;
reg [511:0] golden_data = 512'h0ebbdb2aae4366868c182fdb9c49c632c6d793f197cbc4eeb32253054968e1a86aadfb84fe83965c7da6cca705874f16fe6dd23d136b1fa195ac470f2f4a432c;
endpackage
package dat_24;
integer pat_num = 24;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0aa3120bff64913c6b353e943d4d32066cb5e3064bce750ccae65ad4e3847120033568e2aa13a6f4ee40bf63cb3ff6a42c76491a31c07222c0475fd1bc8fe1573f7e011e5545d39f9be12653b2f34721c70c153232e44c140e47ce68eec450ae;
reg [511:0] golden_data = 512'h1cada0be409961a67da0e929095ecb0330cd463a8834cb28e51e20c0e3fdd002737e5822398b141290b32236fbfdfd04c4c95b6ce02e86ed9b000775003e39b8;
endpackage
package dat_25;
integer pat_num = 25;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2af08f9ba85e72e8b2c53d33ccfb19cc36b6a7b69510ea705cd4d5250e43d076253ac07a6bfbd576785a7a569d2c4322e36da3fc0896e3112325922692cedbfa4a032ff1827124fb8af0d2d60400209437d46c796414ca40fc5f1319da57c646;
reg [511:0] golden_data = 512'h57e8f41bde271dac7769ee0a1f31715425d2be9c887e81f2e240b8984e2a771a3e761048858041d24c8109a77a48bfbc9c39a64616c14a793e938b2200a8e764;
endpackage
package dat_26;
integer pat_num = 26;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0976b7fad2ad436bbaa84e7e5e633d91cd380a4f07a5eaf3c157ae585d521e96672e9c14fda845048f75f2092f64d7ad65845fdaeae4ae4c794eeae0b84b6feb3070ab657cf199af44de9f498edbee1d6037b54aa2638801fddf3fce11241d8b;
reg [511:0] golden_data = 512'h6e9c6633876d5c3cbdddebb07957fdf1f88d97a44f244b24a64f0f1fec67bcc4453eb539d457c071cd8583ebc2a8177772973cefc2641221f137fb8bbf389bcc;
endpackage
package dat_27;
integer pat_num = 27;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h26823cd3a803388e5041856934ae37280104b5b77b1d85124c21a5eefd3c604b21214363644376c0d7c9ae82e7fe1d0eba2817b2cc5e2904f71572651a34da1f713e75222e8a0ff798f4c4d7352db0c00dffbe374a72f32fcab9f5506e10f84a;
reg [511:0] golden_data = 512'h6d4e31c9c156693be8615b9daae992ff8cfafd50ad1fd80eb6b938abf460dfbe68e104a65a5468a4673894946f5b56514f393e9c1dcbe205f19e69295836b638;
endpackage
package dat_28;
integer pat_num = 28;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h45e5d8107104ca598fae636286e237851b1195634a58f8f2936e77ac5aa3f90716dc705846fd7678c1580952590791018acde149b762f7d162a65dafca883d9366d832e326e9455dd844700fa401bbf1cb6232995d25666ba3b5e2526cf464b4;
reg [511:0] golden_data = 512'h3d221c310f82659609c0223e418403bf4b7ed4f2806d95f58997df24bfd6b47c53f9513ec0b9f6f33671c41bc1069529480c2c460d885aa3b08ff302be7933b0;
endpackage
package dat_29;
integer pat_num = 29;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h54eb62aa5d49b2dcfe2f9e31a63ad208d53cda8e47db9aad93e1603b0afc90d32e45fcb02045b8015a6db7904ae1b67fdbdb2e6211f1085ae341a1aed35bc7ac5e2d71a09cea65e513f6f17325d51364de09aa930e65b67edf0aea79beaffdd7;
reg [511:0] golden_data = 512'h0f634d078156cedc6ff1924e5a118af6a75f6268e65da28380c32618556e28f403af1e7ac06893e92a2ce819376d309ca75ee3d46f693fb1ba5e0826795785ca;
endpackage
package dat_30;
integer pat_num = 30;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0ff712816ae5583c9e567e436373efcbc9b144f77c47f17d02fe6830c96ae6bb534453b92068565e69a1054fdfbaa7b9559b8525ba3594feb1db5aa0567073360ca9232999875c4efa4b990e6d4ea527b8106901c6b3110e11bbc837ec58271d;
reg [511:0] golden_data = 512'h6fbc134a36a661cc8ca6f123abd99cb7f3017a709ebd1fcb40a864995c7ee6305484e55dc18df4ce02499d6547c534c8a62c027c85a7abd7240f717af3ddc65c;
endpackage
package dat_31;
integer pat_num = 31;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2e299157a0a2e3c7e399def9175ee8f90f07442217361cf688d2cb7d24776db8000c792cefeead12c1a67410da1e594dba4aec9d0737e5850c8c7c58580e5f38718a780ff6533b5741b728ace06faac38261ce2b6ab68424837ffa547b21c284;
reg [511:0] golden_data = 512'h352fd45d3e14e3ed5a3632475b1a929db6a1aa7a7c8ef8dfe58a287b0d155d0c5a23c68c43cfa79d877bcc9955231913003f6f79bbaa90633a44b52e8c1f12d0;
endpackage
package dat_32;
integer pat_num = 32;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2c989098c72f60745615896a2055e431eab72d477d6a5056863facbf05bb5a615615139f78eb8230074b626c122fcb514cfaca80c346c99ed1a80316c52e4d052c6f0b7491239fdac39c53ccf2319f697c02990c362613e31a15a90938b142b6;
reg [511:0] golden_data = 512'h3d60cc2238f0db5a3071805200170671a0d3cadc7fec9b77a83be351182c35805a0be7abd3d240681f41cd2900eb9ba64135b8887d231ea16cb8642eecd9ee4e;
endpackage
package dat_33;
integer pat_num = 33;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h309ea5339f496a68463ee29dc96a773a9fe20a3547cd650c26a670ca900102d1231ea00533cd65d4a8675e9e5dc4ea6c96020ba3900a2ff625f906cd9695b5320db39e7b872b541f73464c7fc5ce24fb0692c5d3ac8046848824548644644322;
reg [511:0] golden_data = 512'h211feb430c121e20a811afb424919c2154ea9f8d77846107ff507eeb9480f26861e94e01a0ed1cd79d4f632a0a53d7a6a65c29bfc732eabb9ea2545708c768c6;
endpackage
package dat_34;
integer pat_num = 34;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0a582d9c679ab1140869d8f83efa222a76dd6935af157ca9bf9106475b5434230853906ca780404918ad204d06dcfef91e52e4e00de26127e531527cc0432e9d530ea1b8e42d98885b0c070b593a637b38f103a8cec5d7218e3bdd48ee37f19a;
reg [511:0] golden_data = 512'h76a61338777f4cd7ed35f161a4471bc6ed5d860d2d383e71ebc5f14fed259fd0444fa3e676908fc88c929493ac46d3fb616dd20adbe7fc6942848bcf21899f86;
endpackage
package dat_35;
integer pat_num = 35;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3ba84dafd56fedb467b489315703c18f58c759edcaa7ba0ae5aa6654aa015335063ffa5f61f67cf85089dae13e0f62937bf2f0f9d3fb59e284e93b90fc94c5a11e7ee3e61cb67d50f00b6f7afeb8282ffd02d3eaf65bb7d232709cb900b3d9cc;
reg [511:0] golden_data = 512'h772b205bff3811fe6eecc64c3168e817e7c4ac7c9eff46117030a7b55e60490e6419c071c09019b74e1fd4ad022592489879acdbe592406552d744657c368eb2;
endpackage
package dat_36;
integer pat_num = 36;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h12fb816e96c88609caedc18b76da7d044363c364806b11a950545513559e53c864c46b1588fc3488ac81dc6593ccced583a7f0c13762ea7e75c840c2c73935517f26f010c64b40a011da7d42888692d9a3b9e2d0ce46b67a038d179bf27dc520;
reg [511:0] golden_data = 512'h3f8b3b65286ab5b30fff21bc2714427fe7458d062c6cf098a7e7555c2931ce5e3dea273da88a7b7f63a56f821feeb611b8f5efef35af84463eb0ed9a506612ac;
endpackage
package dat_37;
integer pat_num = 37;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7a54439ea71d0fb58bd78a2a2acf5df489801803119f58766a95ab40f883778e1cbf5db880f7a1cba06ffeb992886af01f9e5e95d87911fddb635def98768cce17ec65c83467559f3e9f9e0b1ea45d35eef2d79ab0acaedc728c8b2bd0a11310;
reg [511:0] golden_data = 512'h195b225580b4d3845166a3dcb59af8be0678800563c64042baf62302c4c3c9120b1580ab416ed2ec5e99be3ceb61c990242ab4318af9a29d9e5dd33d5a836490;
endpackage
package dat_38;
integer pat_num = 38;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h583c6364caa84d3d09a8b8cf54d12fa7d42c759e7cd97145688e86b0dad7e63869821310d6716fd9297c1932309bf36af9e7c67c22c8ada178c07b51938de5d046f9085df904a7bf777cb77d43229d2b3c19fbb2aa79b74a73eed902df8cef07;
reg [511:0] golden_data = 512'h21db8c06c2d404e18811b42bec6df1578448afa04f4e0af9ba0677717a2cd0fa31ab70e38c0f1ede1c195e4f2b9083573322b5c35f8d17112698d86f364bfde2;
endpackage
package dat_39;
integer pat_num = 39;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h073eefd75f8e2d8d21b7a4ce0a35b4ccd2b9c5d8892db263fd721d176fe9cd400522626c7af331a27278249b9f66607a6ec390a190ed6e8fb706a3558d8c44666a3295ffb9ac5524f3849e90866833994438e8b7d2bb44d15615ee2d14189b41;
reg [511:0] golden_data = 512'h35735fda7cbec72064791011316297c151f01142edb0db87235af7a3fe7e606c59ddbd30a2f97d9f7de08dd2fe6b6d4f3ab11e35c4233f32fb035f1b8012e7f0;
endpackage
package dat_40;
integer pat_num = 40;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h14dcd38c2f2acade8059d122c44be75e8ec6d508264cf72d0a6fb61456e762001dcd93277a84b083fe2c1cb8534ddf911d6cdc3546ed8d727e29542e69f4b85d326be1f400513669b624db3fd6fa84783523aed9821e144afc5d5f3356b9d1b1;
reg [511:0] golden_data = 512'h4299871d17e1754f31250791f42e8ed62fa2c0f443b6bc3f0b402cc1d2714d961696de1f3ef7939ccd2a1202ebfed669227e03d8779e25f7acd929a634c051be;
endpackage
package dat_41;
integer pat_num = 41;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h616fbf65a96f3a6e328b4a1f7d4c2ad58eefc5f4d1af95425ac80da91c37c34805e2dc3548c688eaf78a2a8bb7444e658ab8ba11b50b54938e6c571267cc42e56eede9eea6607695c470a43df30d70bfa58964869be8266e0e409974aa8111b4;
reg [511:0] golden_data = 512'h4bb864cb2cbc7705e2f0cb95292378f70c220318e423becca36f9b28e8f5070a0cbfcdf0f13808cde129820dcf1adc96289f37d3461f03f072e6267b8f0b0dd4;
endpackage
package dat_42;
integer pat_num = 42;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1ed07effdcbf56a810e683c0fa8af8365fd3033e0c7f53cd0d52ecda9cfaae9b4ef6bfc53cb8262b3b889c916d84821e4554a728ac729c233e65c77b2285c84a1e73fad292eaeaa94d57beedf89e173df7ab5c486914965c14eeeecfd58630c4;
reg [511:0] golden_data = 512'h65526e19e88a5805310b48e2ff6db025a0fed3e9cd88035ba380761e9010dd56235e63f3a2b84260bc0ad60901b4f8c6486c25f31ceffacaee539554f9ecd242;
endpackage
package dat_43;
integer pat_num = 43;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h598ae43fedf55a4b3c99c19ba62ee4355bfd38241a608a693746a2a28dc0eaff1f25c4be815a45d4ba9cac7d201eaa9440221920a3144243d83feda993f473284220ba6188abb5d308f47562328df8a74840d78bee7a426778eeb688a9696b65;
reg [511:0] golden_data = 512'h5ad0e335a4de4e903d4fb4ba61da592ad5246c2f8c928ec28fa4b2a67bba36125ac690ef9223d09da629fa1778c1c77f37b6659082bcbe904727dccbdd887fae;
endpackage
package dat_44;
integer pat_num = 44;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1452e9860fd9561e650ee6959178f8999961380d19367a26d12ab255795fc265524303d987723923d07eb6a2f36f9c436a55c0b580a25528f9a58e4e48db742d2ae98d6159bd7736d92215748b6ee0fbd850be81062015932d14b9fb4016dd75;
reg [511:0] golden_data = 512'h355ef44514599ab0447ebccbea0ab080b26acf16643a7b9bca5df93bfad03f886014c049b20246f0ae72d4f0bb1788dac71366533e858860e49011037ddab5b6;
endpackage
package dat_45;
integer pat_num = 45;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2462109dcb236ce4f01c154e15e9683a1b5b6ace338b82ba7deeac89aa14c6944068a176e3186a5fa9edc9456914e950ccc35fc3089fa6506a83ff9d59d7bf6b5b1b184a64ceba43e20f928e7efe33ffb258ef1676e34d0c7efc4c2a2d432ae3;
reg [511:0] golden_data = 512'h61668941e30a288c780505496f2c08c9f6ccac3f1fd43699df7f91f2ef29b1aa0b375d8581ed1e153305d1ead575ce4b87053140a0085e175d288abd3911f9c8;
endpackage
package dat_46;
integer pat_num = 46;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h47f8b776bc1bfd408da3654df978e27b6b66a8a01e858cebf7049a53db7798380d1eef9ea31de11e20fd43e39ec49bedc7d60aca736044b8fdc54d7c1331b651592e9b4e10d3326b970362376d7623ce5dfee874df7faf052c1fff86023540fd;
reg [511:0] golden_data = 512'h42f6791007b1ba152ba0f410fc5b27a33a420ddaa5be911e03f98d3bdfc1a75a4cdecd681e372bd09b6ae0cd28b74165bd420ac5f89d1329e20c1ee7f25f4a06;
endpackage
package dat_47;
integer pat_num = 47;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h11b895c8d6c7768553aad2fd98f74d13a7825826d697b51d9a4cb9070a10937713d30e21770f78144d233073e958c20abd6e2c7f3deea62c8e08ae9313e4c0a46cdfda8e04fb3df04efd96f29a64f2f6109c569dc61fa4f0dccbbd29c9138b31;
reg [511:0] golden_data = 512'h1fd02ac62ecf56cf8be8b9ac879374e2719e64bf04ce9b622b2e16074b49807669e8d0a369ff4de95a28cbb839a9f9501e46f52a7f44a6b6b300e323c1356f56;
endpackage
package dat_48;
integer pat_num = 48;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6b2aeffd0ab29e9d0129c09926734bbff67536abbd3fe351aa8c32f84b8171bb1320dfe661654e7bdbb1de56164687182ab8c4d146fff30ce1d5e35021daa07e2eb17f440a9e728c18d234aaa068820a758ec8f9c41d9f4057ad28b790b0412a;
reg [511:0] golden_data = 512'h707beb941a868d4cd09d6060697b7c5d4816dc903b3f289191b62a2ae4f6874c29ddb1978d3a05206a94f1ce4b1c9899cfca8115309518d49d66e2337bf71b66;
endpackage
package dat_49;
integer pat_num = 49;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3c0929026da0cb7d172c043ba5040d0c66c6773c20e6006a4eec5187f264815b2b793be9307f028b7b66ae1e6f35856f89f0ce17cb12d3cd272e1734af98f8ce0febe3b96ca80c1f76112aa5d2eaded05c49643aa1a8bde3d46eb1ac608a9967;
reg [511:0] golden_data = 512'h7577d6ac852c4054d222266bad745ecc7f59f3566c0527a305ece762b37805c27f82e1fbe5ce25c0badee092e5407a195b34b317a85427a1ce7ed8109390f23e;
endpackage
package dat_50;
integer pat_num = 50;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h41078646f523bab911e4ccbe5b93236a2db666beb617e53f3d1f051cf785acb93ca002cdae31eecdaf5a835b83847d1f4947a8aaab1d701a8141a38fff2987464a4229704188cf4640d1000ec1db3cf17ea7a366f0c0a350c973515269d7d2b8;
reg [511:0] golden_data = 512'h398f8a8ea7fb6f927b16c6b03df132e493f7fc78b5599770819e07ed52ca8c1e69336d5d30d4443e7bc3dd4fa8b1205629f98f043a6ac4797d93649f6e1aaba6;
endpackage
package dat_51;
integer pat_num = 51;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7e44a505c6c2731c69d367fc0cfcbff568f7ab7bfd04b8c29aff2d955d1d1a9412479bf55fb260bc7596d7959c09b95403b3296c2ad106e74505b50ea7107f5c12cce817ec855b5abaedd80e8ad767a5cf6a8c4c1b88196472655b412ee961ce;
reg [511:0] golden_data = 512'h5c4b207b2eafbb229b2b556eed3e9e92e520debdff34f819c191b41a96fa6e0029d8da25317c90cd4a4a7fcf92c8bee6f8baa5702bc5ecf2763b7815bbf33672;
endpackage
package dat_52;
integer pat_num = 52;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h505360492a9c759fb53c569d8a1ebeb805d7a0162f95fe630fa049a62ad8986c4d621075c1c75edd40d713948e929a55f387278f0d9b29d50dda0eca96245ec007992ce819a950c29e42195d5d0a6a6e67cb614bd7bd97b9252c212f1eba806f;
reg [511:0] golden_data = 512'h1d2f17f45118018de44a575c8052bd6340c530b6cec4426d65afa913b8367f9629b19683ca39ab598e13e080bd89acc12e6ad98f978cddf0b42bdc3aa3cadb7e;
endpackage
package dat_53;
integer pat_num = 53;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4f9a80d373890b7c7145d1908a397f52d3856666c8b121322484cb83b9159f1b631c441c77b2ef2cf4402e500883e581de1c50e71dd1b053fff51e9581bdfada42fec33339906ce22f1accd3166417f32dd51c5d7d76d038490fd0c2dd37685e;
reg [511:0] golden_data = 512'h0955c6c6de156eb4882a980af80e0237476edb4d9879c0a85e2ee5f5722b604003a8116e8224163aaf0c96a80c1d9b7453d7878f36dd115324d914c52295af14;
endpackage
package dat_54;
integer pat_num = 54;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h77f6cfcc603f10d1abd6b895fc45301787f1da922259fd0128bf21cb800cda1b30d09ba4e9da30579b577b1e57bec17bba1ca71d4387c09a275a1854d05fc7277ab3de3e7440f4573c373504a7ac5828c323ad29ec50b364a955a6dbb9d0e7a7;
reg [511:0] golden_data = 512'h239fe045ea245fb96b2e1f3f68ed793c33e387f32e3107e5f9e18987667f6fae4fdc302b804f80b0964340f38c81db8a8f82525b51d2663e96a30011c205dbde;
endpackage
package dat_55;
integer pat_num = 55;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6ddf88a978042752ca2b10bc2a2775d5e1d0ac69c90a98047a0e6f69d1d763fe7f742074979c561d0fba6448cd29a9f128d0b49ccca7cc7e0de27aaaf5c7cb2c5a81e9be3f3685e9b930930d984f2f2344336b13737c15a5ec2d9981a4f1f0ca;
reg [511:0] golden_data = 512'h09a6e0dd1dc8c66638015514a802ba5f68968966d2685baa41bc763d63c9c2643c387580344c5d46cd824c155ee69c29b7a3cb637b55153f943aeacef2be949a;
endpackage
package dat_56;
integer pat_num = 56;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h70c1c00eea74a79b5c8546636a45a2d23550aa820fdd56f82fd4a5d335b857027d2b0428b16b190806bf12bda338ed7e63dd63ac8e295850a041caa49cf5079b369506b2d225e414e1e67c7f19049e3fce288d148adb75e6b3ba1f3f26a69447;
reg [511:0] golden_data = 512'h1aff380b686127dc36a5366a2d8d396b0e9f25b1bf5a447ab43e59f7ba3ab70a7223d2757cdc8005d96040962bfde28a29df7abe368851f46553de49dbae0ad0;
endpackage
package dat_57;
integer pat_num = 57;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1c52db88ff9340ee564477ab2b970ec4eaa7537166d1b0ec5e22219c28f36c6826b264023f2dbb0008294e563bd375cd8514e851231d9b06d9b31f05baa09fb87579c567157898c6574aca7a7ba85228eeed5741cdb5d77c85c957530a7c625a;
reg [511:0] golden_data = 512'h5dd51ab7ad0eb725e5059c54c14bac595fc82d017f5baeae704815dc2c25fa5e363e66d95217b83203185a0918d5a8aaebe7a23cbc3188cef54ee897989232ca;
endpackage
package dat_58;
integer pat_num = 58;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0752ba40d1f259b704ba11b5e39ab8a9aab27f238b32c8a0f7fbc1df919b1efd418dbde7ce1aba881783a189e85e6c93759bbba8211c8362e0d3a2de291549a4451bca61243fce214fecbdee63b9de3d158921fe541db23b5d37c5064ce46c87;
reg [511:0] golden_data = 512'h233fdf5cf3ef63ef264d062f7ba5dea4479fa65ac26a64332918472bde30b2be6e620777d032379a3260b550bf8e632c87446bd8fbc32c3741ed9922c000f0d2;
endpackage
package dat_59;
integer pat_num = 59;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4ffada53f6a29f5b0a1d9b52ac41fb004740645af1e49e9b17c6b988a63a9fe116f90fb4bae224b0c3017018917f49dc49f985663c93d571ac6bafa157d9e10c01a8b5c1167555cde981f77e2ce34113c1b0d884b30d0b449cabc87bf4688dfb;
reg [511:0] golden_data = 512'h240bd1d4320a22028110c77935d3b7818881d6487cb4ce4541bfcc22599a56782c4f6f6b0b3fa2b1ddf07519d53011e16040ea7552863fe5a2c2400cd2d9c3ce;
endpackage
package dat_60;
integer pat_num = 60;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6a788a72a0c92279b363c2e7744c0e9c1c1b5b44349b2b5b91d8987f7cff84ca3f18b67289927ab86af418b9f8ba7f6fea648d313a7e4580c109fb4dcdc72550157abe5883a8279ac94f7ffefbd3e286813dce9252a201429df6d8ee0af3491f;
reg [511:0] golden_data = 512'h233cc4491cf84276599ace045e368bd90b642d679c477520783d7d6052e875fc3d97dc1b22ff7dd335ada39ebea500d9d9dd0705878b00ea444c2c1af6ff5fe0;
endpackage
package dat_61;
integer pat_num = 61;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0d294e8411be41314d29bee6451be07bb0b0e45b4a2d61d98e9ab3571ba7a0ef2d977cd5c0dbc8f9edea8bc681bfe1e1f8648c0d231f8d193d964ec9577835471b1e2de1fccbf920536fed64d4cef8d9dcfbb259d064550b1541ac3489a005e8;
reg [511:0] golden_data = 512'h5eb9326e4624f691374eba75b59168cd07446aab373ddc1fdefe43a47a5916da7a4faa577edd9c86be53abbd795158ad4cdac8f97dbd305f88ad93b8af3e6958;
endpackage
package dat_62;
integer pat_num = 62;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h04d0213930230a4fee033787505b6b38583e60d8e1cc2c482c295d45a24839347f77c835dc46a44b11f1fea0c941472fdf6ecb4146a9498d64129228518484ec4e5dfe3a48e0faab12841ea3fbc49a1bf93a9bcac32ba7d2159456e66f9d3dd9;
reg [511:0] golden_data = 512'h4d0b280b108037162a6a481bb263f7b30478d3d9bf5755036aa49bc173e3f37679aa3c39be05529151107dfdfb009af8dbbf1da43aae5d79aef37bf2bb68b982;
endpackage
package dat_63;
integer pat_num = 63;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7f2d09614994a3b899bf3eea93221d8b154048d5bf2498e653b75fc1cccded4a4d75347daca713a54c05399c27700b1793cae340b01fd4f707b5d08321808bfe366ac07446952948db961a100f9812a1f32926fca2207dad985c37307735c3e9;
reg [511:0] golden_data = 512'h786c3f9c9a4ea16493b5878187986fe548c280ec2131f5b428fce5882fe644f869aa29ecc7992cc376fe9e814f469c6c17f3e43284a074c8429c4594617b8252;
endpackage
package dat_64;
integer pat_num = 64;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h30b14c7beffb12f24dfcfab730a3e80401e125ebbeced108fa7fe0c48d11439c1e1fa235fd4872a80f9e9418cb8fdd1037ff1c4b7c4a625ce779da56c22429097ce22a47a540124558b835db43c66a80546c2c7208a64ef440b6e3c0c3958036;
reg [511:0] golden_data = 512'h05b723a73b66eb2292ec8e50461590431dc2d5bfef08f335b4af02b29d5f912257c3e98aa385f3797a2fc3101a533f8f6bfae4fd2b6ac8c16c2514fc4594f79a;
endpackage
package dat_65;
integer pat_num = 65;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h32ae20b63a124b1aa4a0f57a9a59f5e66df72523b460476111b2955bfe3ba072753dc5fd047f6c1be997d6af76747460fff502b921b7d973d7b5a490fa320ffd1c396bb473ca377bde59c9874f566f40ba38dd8fc5710f7b2849c4f1a2cc2154;
reg [511:0] golden_data = 512'h723f60a8d7bed7bd2fbffcd00d357de3584cc0ccf65e59f1068ec5f0ebc87d462792a3bbecf2d27cce55c6d672e4b8c0fabfe461528abd14cea90460932a0d74;
endpackage
package dat_66;
integer pat_num = 66;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1e941916b19a30523f94eb08a89a003758303bf7be123c8e9de0a95f29651e7e7287235fab11f804cf4227790876933c8784310d170a6cee92cb710c3c04db6c24f59ac340b2229c4e3ec57d5942aa34fb7a0ebaa6f6c491218350bb564afb27;
reg [511:0] golden_data = 512'h22afb69151809fa54aa711b991785446eab6b84d38a153adcf9bf537a4adc36415bac86f4fb41d42b0294686f158c4cb24036ce6866d1a4e787098db5d4b0634;
endpackage
package dat_67;
integer pat_num = 67;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1017d9df12cfef367686a4640179c9f4d45880eda44fe87fd96df9f65a1eeac70ee2d3e68a244d07b9c10881c04900efdbfea9d74ff12720eed448d2d6a4d8fb161ea5e892c854c6fbc2d8c1544dbb54a9fde65f8c3e655a6fe3c341dd48bfc9;
reg [511:0] golden_data = 512'h69a07319ec236710b010212dbfc2e187450388a23f2edf363b63780df71f8c583606d6f2020c3106538e4a6b0d76b16f732bb7d316d51786e063ef873d304fd8;
endpackage
package dat_68;
integer pat_num = 68;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3ab94d37e320ba3220ac616fa19d8a8eb41bb12a475c8349ba6a491c4516126b626c15547c4cf510a78018d71560a45aeec9b60d10288d713d7415d7a4c237ba6d1f7c43c9c06bb62eb1d4ec4e93106fec559c6d660cd75818766215b47d14cc;
reg [511:0] golden_data = 512'h56ebb2ff20ce922925a211e9057b4f1732f5c5c699b67e873d0633d1ca5bb57a63c03df1f8a25f75fc2e5a11fe09486fc5ed6431a04fff1b2a114f3d37e724f6;
endpackage
package dat_69;
integer pat_num = 69;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2473907b3657f732458ebdb48b43905c05a29180e58a47e289ec00f33a1a5d2e2de2bf792534bf4202990256f55fbf63761f31f77f76a9b30e19acd470437ae40813224e20aff57255ec24b66d6401b32f654e38d6c1f2ef783ec6e5ac0e3c0c;
reg [511:0] golden_data = 512'h5fb445bd153ca5f4b8022ad48871b151b683bce6cb9651914ab7e591fea4ddb8481ebebdc3a91e6d4eb036f9981793b100012835e466bc90c30b6ed9b6064406;
endpackage
package dat_70;
integer pat_num = 70;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4a4f41bcbb8de61270c34f887d284ccb534ba9e433d2e46d4b6ab49d8b331cf64a4959616633f9c0d7debf240e69915e32539eb8145600893868d461e0fa8d4f280d3888b2def5c7b4a214cca669e5bcc9c84160a219852c389eb0e17bf90e9f;
reg [511:0] golden_data = 512'h3f40dc59d89bc74db59397d1be41ce1004ad185b7a053260eeefda9bd36a68ba2c6b256bbf0187fb8e03fb2b9e83fadda2c6ddcbd3fdac257ca7a1ff638775ac;
endpackage
package dat_71;
integer pat_num = 71;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h60d94aad84e068055bcc08ed4533dbe23561070fc596ea4aa899e1fa538495f8485cf5dc0e87b2b8d4330cd264644ce12a4dc77ec57b5c325406b12682919e3a74cb1ae589bd692271132bb7acd2165b266dc6015a3ee4f17d949a661a933d96;
reg [511:0] golden_data = 512'h53ee04597cee760aba3deac0aeb37222e656883e77696811826df6ca33c3ea5e699f3c30abb0f2e03852fc66ceccd31885c0d8ed281c810400144905054fc1c0;
endpackage
package dat_72;
integer pat_num = 72;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h05198cda112cbb41700066b2b1421f5060a04d05508620b586f8943e53d4a230615b6ba9e0db4325e94ebed8d68c127951e77fb3713114b05a9d682e229dce4778d880436a87d01adb528a849a059e8ad7f239f098d648996692f04132d126bf;
reg [511:0] golden_data = 512'h4fa23171e6bc330b90ec3c5351f1c3ab2683c20b1acdd7d3d3602445cdd93f08591b1fad36e256a08f5b9922f6edcc5177a20ec3fa3e1d4694b2cc7ef79f7b4c;
endpackage
package dat_73;
integer pat_num = 73;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2418ffd83d55423ec808d645eb3656539076932092be19105db7434a36ae05574f327f551b9b8cecf7541d9a05fde87b1b9eef95fa290bdc3be4e327f3a1cbba6cbbbfbce94a17cd9d257107c799639e7cdf293700bfefcf7602a566e88446d5;
reg [511:0] golden_data = 512'h6ff97ae6c3da9d564c3c0315f1a74257f0a873c67240c33ef5575d60c8c6b5162fa980f59a6b9ed8dbca466519c9b2854053cc9cc40aaea5e6e84af229780bd6;
endpackage
package dat_74;
integer pat_num = 74;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h29fe241e778b39f165a7fb463491adde0f85d4fccaa9a783013a992f2f1081a16acb730eaf0ee1a8287a205239278d91a43fd43b1acf159c4635fabe9eb2c8543ca7cfc9f9b0ff7dddae42c146d5144a60a2a554201b366124cd18d3084a86bb;
reg [511:0] golden_data = 512'h0c6904c52d90c4a3909e70e22f22df4c4dca4fc88cc7abee03d3076fe420c5fe5708806b396d81fe764a80beaed74f86a63560fd27c3ec88b94da1ecf7fefc46;
endpackage
package dat_75;
integer pat_num = 75;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h08ce0d9110b173bd913466c34a3413c9b2bbe53dbd74284cf2f57b53be4e1adb38b95c04d8b1e144dcc911f31ee890e69008a6bd38ea377dccb8093e1704fee802f5a52563a0a42984ca7cf1f5b4271e43b5d4424aa57e18a0159132de79f899;
reg [511:0] golden_data = 512'h6326fa15190a7f81241afaefd1de82c41f366718b086fbf95de3e8a2f1675a682c67091153f6c92eb5920811692426c28a75e5a7fe7cc52d29789cc94cadbeda;
endpackage
package dat_76;
integer pat_num = 76;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h605b78b351f6547df081735dc8c9fb151431ac930ec004883c738d52004b5bd27468531e5fcba703c428954f2b57b48278fb2d14de0aa830d249736f4bc447372517824b9419f4c0d6155cc2327d8727f9d58cfe4213773b495b2e6e24982e2f;
reg [511:0] golden_data = 512'h0c58b3a4802e61f40ed00d4c88f43bcdd20c58c54510c1ee69f7c11bb4505c6266fb3c5f6a82f27b90dbe5a10fc13a0f873ef5913c9bda2de0ee3b9b54742ad0;
endpackage
package dat_77;
integer pat_num = 77;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0373eb62e3adbfb1a01d24a0f0a59cd6e17877cbcc1257a0b0d1ea789b2ffa3554db3416c63ab3dada98b3edf66aecf403d9e78294ed0c1081b35c65844b744e6dfe874c6605fee59fc63228970e797bd090364d9322ace840cbf66a1887562a;
reg [511:0] golden_data = 512'h5492293bdb4e2a03260ff33b6bf44dad509793dd96e46e40cb6f12c6ab2a4e7a3b6aee48280a29132c00c0d5f5c994e40c8fdb118f92642cd91c2621296d3eb6;
endpackage
package dat_78;
integer pat_num = 78;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h11ceb4619ffb751339ac85de7deea42650998e7cd63fbfbe2573936004f8db284d6e08bcbae5a0e1e71b2d9e3a9732d584f3c4ffe9a24b713a57762a5063b04361f83f4c7bbd3d884eaf9aaec2840a30e4247f15db287eae2ddc064ce586c6e9;
reg [511:0] golden_data = 512'h37264e0d8d04fcbfac4a342aab1ee10d7310a337a06c0660f956b29114f8f2c82e0594eb43ea5d272954942c3d8ace9b8d16009f050aeca17bd64939ce1b2614;
endpackage
package dat_79;
integer pat_num = 79;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7d5979a0f95d6b3fd04ac37820470d7ab2206dcaf7c600fc79e0671ebd2e803d736f8039a339a8f6fd7b4ba19b0d509e5a17d9a28fac9d01d85a6d4aaa53f80e26972e338d732762afe05828aac2935c583c6d96876be49b7ebbb714af09947f;
reg [511:0] golden_data = 512'h7cbb19891310e0f5b7288f5cfd795600db72b7251a9f74a2ecf2c6e02ac91a0e03d5cd817c570152d5ed4e23512ca49cadc1b856f26f5c569debd6ea8f4206ce;
endpackage
package dat_80;
integer pat_num = 80;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0c82852547d608eb1d1fa9a816302ccc90d486c1f305ccaec1e61283f0f42d72504462c06c40ccf6b52c49bcad888288125eb905b83b38429b1f1ae3086010f562665288d655f9deb780dd671e16e55b7f87c99bb390187f9c0d61411d284cef;
reg [511:0] golden_data = 512'h265ea06b23abdde3da125fbf5a2b095d4f7b88c62981758f02206e2a8b59fcf061743f3ae878af3c5e93214439b29d16c9ac51bfbf8f9040d2b27ce31c66b6fc;
endpackage
package dat_81;
integer pat_num = 81;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6ba610bed0aa840ef63e3d85963ea93e062e80a559bde618e77a39e2dc2b8d54286f78c258f7202d81d35255f3ba9e91f23cdc5b7878733b3d0c80a234faa59947175809c071e07d83c3b6bebd52a1173d05ab1ea4963893d92203f876ca037c;
reg [511:0] golden_data = 512'h65f05313beb5b5c06a3a5f2848f9c59d5f73a4d54a8380c0da8a2e8b7c7e254c161e6b174642e3135a5d553ce597d351bd7dc84618b3fe507e6d8cbbe30cea9c;
endpackage
package dat_82;
integer pat_num = 82;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0a76d745692df277839de700440852ff29c8b2694e7db2c90cc338bcd3c7c93969134f0742729570d733743e119a82559664968f5306c62087afb0f184788dff516e078b0cff617edb348568dabc76d6584eac98602332a062760dc5211fe23d;
reg [511:0] golden_data = 512'h50d8d54ec8dd2910d2d122c0f4c5ebc37ed7f516659d3698769ee652abf9ad8871b37cf426e30c0de5e4e7a2fddd2483afd2ef43dcdd9f530923944b248523c8;
endpackage
package dat_83;
integer pat_num = 83;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5339b1e68459f58d5c3b6db5ff968494e8ba902c66aecb437d8b4ad17a1136aa48ec726e91a4c0ac8a1889179e5deb7e898d297376a15f8f4c0d6834694464b44a2b7ae904038fc7df0e02140677cdb135a41373dbf8cbc0244702a5a2abb3ea;
reg [511:0] golden_data = 512'h511477ba207f9fa2aecfe189fec6862b762b21723bd39ff380a88242cdf94b6e50d473a8c64156c0ae37dfdb7de21bdb7ad5c70320eb4dfda3d481f1cd588c44;
endpackage
package dat_84;
integer pat_num = 84;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h65dbbf5a2a45ee9ffef2a868f7ce0007d6cd65a55d3381c4a4efb236c3d931a955121ca41c56efe16f5ad3bae1050b05ee2ee98cdbc93b9c5c2374b59e8ec59c72e5c9a2602d8bf9324a554c9a81db248a3fb054950b9436cafdb64f7c4024db;
reg [511:0] golden_data = 512'h1b6e1d1e2939a00d76d9c14c70c0c8acd32a9903de57763956dd6e472978a7ca510e8739fed8c74e6074b5afc2904e36a64cf85afc0ff931289a3f247ec95df2;
endpackage
package dat_85;
integer pat_num = 85;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2447ac7d93a1d0e52dea55ad2f1e56c25cd57f1d1b1f1ea6825f674f6f8265ed1a1d974a8e8e912f9fd5b204517c57571c19a3e282df1f7141f1a857edabc5b92d4e14332a8e0a10b66f488ee611f163fb22a8c0d3dc2c5ea7d005fd6de6f48f;
reg [511:0] golden_data = 512'h1afe3e840dae42a751ade1987bc597dd113ce952eb9441200fa11173da605fd60d1b2e7d153db6a3bb6ffe4feeb82dbbb8051a56c43d4dfc3277601edd7ef2ee;
endpackage
package dat_86;
integer pat_num = 86;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h255bd2b1aec14f1863a87322f4f7c88a47547ab8c646259d901b82435a2159f327f690a7169cce2ac628e3e539ee1ac5f95604ca4b750ca8a76bbccb8fba95e972793920abbcd4cbb7e1d10450c19258e723ed5458e513be8cdb758c81ef3b20;
reg [511:0] golden_data = 512'h70e6ddbdb0424421cf63adb005d2b6760bab0c451695201882f6ddb3a27efcba36777c4861b35c60cd30e10b80c52b221412b16849e3a4367fb0a131ef0acc90;
endpackage
package dat_87;
integer pat_num = 87;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5e897d97f8a068c64d754679ed6353bf224bc62de847e5cc1c9cdf8700af9b7377c86091df2786c641998057e8aa781932d3b5d4a67fe442371f1840a55ffd8436477846186d6bf2a86e93487caae85acdb7d84d2d5aa05eadaec664a729e609;
reg [511:0] golden_data = 512'h7d0098151ff3b03233e75ad4e45797c2c6ec24180f9ea4f46f1eb010299e56b84788fdc67adcd7e0563b3fd943336557d6a43a3312e0aa9e1be2478cb3370508;
endpackage
package dat_88;
integer pat_num = 88;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4ca7e3ec334d172cbc444873a1d13d91f3b47d82c785162a96fc188b96a0083e5c331090914f1f15ca68f34dbf96e316ff05c552ed4e6d519cbbf604dd170b1f43b797699729cb5448c682bb1235c98d0f3cf1d7e9cb3c6f80c0c82b68714eb6;
reg [511:0] golden_data = 512'h57e0ca91ba7f17178df76fc997261c6bbad1d657d52efb7929f2df0811e9de5e588ef353244d8f42297584c7aa5cf6dacda663d6e25d6735e9f616aa73d576fe;
endpackage
package dat_89;
integer pat_num = 89;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7dd62b0edff7df1733b8ebcf95b4dcea21fdb62b64bded526821a1fa44c215be3807a39b0c5927b9d60a6336f7462f606aff68fc9b4b8846de484f1bdd8b3709466634cedc19c850041c17cd50c145fb171036b66c3cbcc1fdbeb430048f27ac;
reg [511:0] golden_data = 512'h02fd8fa770823c8b8508c68e57df1965685b461ce31a81b2d3b867221fbff31278669b624d45f81a45ecbd31f41f4b4620b6fab0ca2c61d57e3bda7bf9970d76;
endpackage
package dat_90;
integer pat_num = 90;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h50e6d413056748b7720f690bb079031cba5363c5630793a8110a58cb43f4c49c223da5f5a7f43bf47255d51c262b486e9e82c683fea6e160b96261997c9dd00d3d5f8ee512415cd05ba80bc877a27194aecbf0f8e7932deba0333a534a89fbb9;
reg [511:0] golden_data = 512'h48d3a75add279129ace64b6032bc4d3e60f0908813d2edb22058502594edbf9e1d37831930475d11c91513347a229e6dcd77df2aa85fe34fc2c399ad6c8260f8;
endpackage
package dat_91;
integer pat_num = 91;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h41ff0d4d7c77a75ed2a905637be166e167673195055e3afe111704a4b9337bd221d540a4a94cdd8eaae4ac98a94be2d1e80838bea7c4438a13dc351fceef482b3cd9d82f9dbacb505667716e5382f7f7ce4efb32b35546e061f0db42da821552;
reg [511:0] golden_data = 512'h0ebc537ec23307b0b98cf3539c9bb5e2c1a782800905fc64ffdacfbed2e57ff464317635015c473a37b3cfe204231a2059f85a1f7fdf3205def47e524fcc111e;
endpackage
package dat_92;
integer pat_num = 92;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h79077f5f87b791bf717e48735bac114020735a0f275719b29f0ceb089f911e7669fdca444d42b392bc1ebd55830dbe21f948ec9df43c3070b2645a2a8aa46822168553a597a973e5ac2f5364951399161ae4a4450551c09f647ad7391f2a5724;
reg [511:0] golden_data = 512'h183ce7d5dd2aee594bce6bb2cb7e4b777b59b6102e98f178efc07013f30563302bbf197f6a5508d460f69e9e6dcd0b529852fbbb6323aeae408eac58788cc3a6;
endpackage
package dat_93;
integer pat_num = 93;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h34f9bfe9bcf5c5e6523fdf8f523f793cfbed1853d35bedea5dc502d594a993b94689f2c0e3bb6cb58864118ba3bef3438a3bbce255b26b2d0c0a0972877f0480102bfce344a96448864dafbffc0e0fb3a66335a738745ab3b5db22b015822e12;
reg [511:0] golden_data = 512'h39c61731bcd568ed921ee1d00cdabfb695e221fe7aad8624e44a2868a369cefc2d2b999b37bb0693490f6cab8d9a70ed92dc2d7b547f7769bb35db444b28c1a2;
endpackage
package dat_94;
integer pat_num = 94;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4d7a5dbc4c26d9b701e01068c1b531b2e59ba37f24db0e900a3622861f60716832de2155933d1dbb3cbbc3cc5c45837147211f49b462464c9fb8f5c030dd33960b30d22bfe9c9a73dde4e7ca15d4f999a4cb283748c2ebad64a93ffaa0916491;
reg [511:0] golden_data = 512'h1930c942df14c9c74185d0f32aa3168fccd1ff5e9d73dda2ec398944cae97c22329ccd74a80cb52c5fec545c055ec341f0f0870a97f2f7d713dacd0837295822;
endpackage
package dat_95;
integer pat_num = 95;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3c0f6d8d86b46524eb91251ecd64139de252b7c6b3142cfa4e06dba2880a37d832fffdf70ec2f2bd5ed39681dad15ba7a2b94ee2fbedd97975370da61c0d4a5f0400f03e438dfde270325e303f09ae13a191263cd06067d145eb5f23eacdef65;
reg [511:0] golden_data = 512'h55db5609d9e7f0a849c196c1740e5b24e19a9d12f15e36b50a85e721e1125812288bb0b58207881054f614762306a42916b1e7388242df29c8cc7463b46a8b78;
endpackage
package dat_96;
integer pat_num = 96;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h09b9f833c413ff69506ff9878ced572fd61319d49e4acf8f1de591038ad290d31c6da47c3190b001a622eec7fc8d3b798910e225cf9348eed94fa741785b39d57950c77cdd4dd4cdd8102c65ac8f84536e44a476603697e755bcf6751ff6c1c8;
reg [511:0] golden_data = 512'h071eef838accd271f62abb46981abf2b7d419f016004370b22992d4db1675c5a7d51fe57415d588d9143b7d13637a840a5ab82d9e70a473e6e06ec765e7e02f8;
endpackage
package dat_97;
integer pat_num = 97;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h69f75dc3fd6a6e9e698382ef68b87ece57b16b6ab7266f3d00ff34502f47b9e4228a6e6810eee74041cc542fb4c93a7693bcf0fd49d5bc52bee31c19bad333ea493835f4359106940202130dc76eb23bdf11e1400c0171cd12226198242c4cf7;
reg [511:0] golden_data = 512'h0fcabe9b7c120a2de8b4c9b536afed5912c1899d704b3d6718507b4d976013b47f3d305d1f0352de3b342cec1923f34c30d8e18083f76575bc3e58d6caa40c8a;
endpackage
package dat_98;
integer pat_num = 98;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h30959f0f3f3dcd53e50b75d2599feb49ce714000619bc86baa15dbe42d760b205be9fe59d6c448918c404209e51632e1527a805614aec22d003f42def9fff0e60874a038f137e81bfee1c99edf1d7311dc09d9e6428c3a8d490ce7969fbaab58;
reg [511:0] golden_data = 512'h209a7d1be4c991f7a02725371df50d2ccd86ff3e61cfbff5a983cff41b99aeb07d396e4c5cf3457c69955e29be74bf78ddef514e0a6129c12dfdf65ccbba00ec;
endpackage
package dat_99;
integer pat_num = 99;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h78c8a82905b0b5a8f097c3d74a2939c4316e0c7bb2fba5ae833f6ba01f16f0667e0d47b515e33306228d3bab903b48e9022012d2f5f461bfd36757ff1a186da1525bf679cb69f67e8ba11676ac86a8c1f7c189401a5ef93d14ac90a711bdb233;
reg [511:0] golden_data = 512'h519a351f2e778fbf2f5539649cae474b1780fe962a334c7635eb873225638b8c070e7c78d7323bc982a5399c3be38b260956af5983e7e93b50794c655090f3be;
endpackage
package dat_100;
integer pat_num = 100;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h02d2cd3952d1843af0374d59be208ae98821cee70ec2c04111cf2862f497a45c34049b5eefd634aeb00b49edd0277b255f8cbe23fccdeab90dba10bd56c5166a00f2faac92aef98182e35428dac1806e3a79884d125dcee3cf2fa7253ce14769;
reg [511:0] golden_data = 512'h0dc66119400d296b5669867b9d0289f1e3f3c5eef93d8847fa373da79042bf3e3c772871d50fe1c5368931c4f587395ee6f28d15f9960ad5c25a7ab995a2fc86;
endpackage
package dat_101;
integer pat_num = 101;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6b47c635f606375e5b79473ae84b9ba3e93d6ac3cedd0bc6542b9ae2509e88f50279c426633e82e8bd92b5d9c792d63c9eca3955b6c1c7c71f63550972bf87105f2eb01baf5afbbbfd615b5f5253b1e7be93b0b44738dab19a0992fa2fcf8f2d;
reg [511:0] golden_data = 512'h4905b725c79f5a57587baeeedb23df21d660966d618ae555de1b484f547e33c06fd50f3a3908826a769045c61acd5cb63fb2ee7e0094fcbe6fb51bf588cd7760;
endpackage
package dat_102;
integer pat_num = 102;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5f2642b43143ee6672be0164a32f2131bffabb56d2b40c47c1b33f450595a14436f3ccb88c5a430ce2b98b371bbc0c49bab6c35e0c5716a057f8536b6937ec8e56cb3a51f1963054a83a06a9560a18d55ad6fe5c7218eb8db9e3f3e5db2dbec9;
reg [511:0] golden_data = 512'h1be13f45452a46d76f7f2dbc8adc82eb28ec5cb0b4d5b6a1069e29cfa87e021a276fc14586991143af25550404fae62235367b1c27fdf5aed3ef1851ea9b2722;
endpackage
package dat_103;
integer pat_num = 103;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3aded0dcb722d896ec03bbdbc47c2a27679947e7e7e5c422dcc2aac2da18e8e92306e22a71b69f0475c8c616e1d7e011b65b1dbc1b1a6708eedb9b78765971a33038b6b6fb3dcc3a39077b45a335f81354d16d172fd14bf0c4b9945911470e50;
reg [511:0] golden_data = 512'h2a8f4b1ff49faf4e790b840f012dca9ea49fcca6b79987ba89af6e5dab44623206b75e22f57ff55a55a1985569d92c25c33d5175329adb573d1e49bf9a90eb90;
endpackage
package dat_104;
integer pat_num = 104;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h35655a18ae97c121a358beeb5e40e7d9b9c1cc86e1a1e2bd870baf5b3d90ca962356925bd7bd2674cb09302367ea4afa0d8099db6c32fe1eda4815f5b8fd180d757d1d651c4460932265b9594f9329629069aabb2ff922c1428d432863d06eac;
reg [511:0] golden_data = 512'h415e0789dcbbe12bee9b3a9206f32e25c2ac3916803c69bc699718836064014e1d1c77b2b7638d94b0da596402d8ba82105b9fa3d21d4086ad681a785fff94e0;
endpackage
package dat_105;
integer pat_num = 105;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h271815fd33d703e5cf2f9227f136389c43b98a7192033a7715318b701f24bbce6734bb979fd4857c39422fa0f4f3c3db5a2b6181e9af7ea3de598216aa7b6bc76320d9bd7c4f53b47e1ca84b83096996aff819cd5aa072f061d0cb3222238bab;
reg [511:0] golden_data = 512'h478e884dfa6c495bcbb8d822b726896a80eaf724a209be39ba755f37f48f42207b2d1b839f6ac3855583cad8d5653fec5802db388838f872a98d4aedbf6b64aa;
endpackage
package dat_106;
integer pat_num = 106;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6d88ac8fd178f65b16707b41923ddde944c4657eaf55204d27a51ba225f6a45438fbeb0c6b77f236ce6c662ee0aa7bca93eb67955d95808cec74a6e93698c52934fd36bb7ce99eb236becbc90281af12ac969a01c2b7befcaf0125b303edba55;
reg [511:0] golden_data = 512'h555e8ce03749692cfe6602e5009f3164ee125bdc4e0d8e20f71ac4ff7357ccce3e2111633963bd8e1edfad03ddc2031da821fa949d6fe299ae2fbd21c3b2c93c;
endpackage
package dat_107;
integer pat_num = 107;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h246cd5bf2656f1128321414995a20fd4b940a866106935438b8a296adfdbeab13bef571aaedffe452c059e2b790600830fca5bdc14b626019016b4d88e2032185c76ce94a5fec5dd393dd365dc8b7d8f90f311318b6e2d88b85a749f2c0f80cc;
reg [511:0] golden_data = 512'h0b9f56601c6456d2ffef3291706c5f5d75fca9ef046553f45314511b00dea1da0f6bc211c91262c0527a21eb2c3b6533d2c2481fcf631859f0413853d3b448ea;
endpackage
package dat_108;
integer pat_num = 108;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h67f3c042b32cd844204d4477e2fa1b980a9a3c9e5075c9926f242c1e0b77bbf32f5401e4d189ac954e6ba48f2342855e7345ad3f17e92cf0d77b74c303558ec27fcba8ea4bd9f3d667279201cdd91a9127d1280e70b36d86dabd6ec00bcc9d2a;
reg [511:0] golden_data = 512'h25b4dd83f7739a2236d24de12de5b3843b5cabe8ed36bfeb773016cd80550e8253bfbbf98ded475a62d47d9f9cd94e28a5afbd4e82be207dfde187b7b82f0e4a;
endpackage
package dat_109;
integer pat_num = 109;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2a10b35dc0008690f5961c76448a9ec685b6637bb2bb33e64a75a1bdb23bb3677ea1656aaa4c65c35b461f2aa7918f7d533632f9cc64b91855b628ff1e883e2e646fec6de475a7b98ec7124020891ed7002b6c605a7d6e626aec8b732f5b3a8a;
reg [511:0] golden_data = 512'h16139d168417b491c67f166ac94bc37e6ff9fa55d00fecf3ae4b0a6a0541ee7052f6cbae36222ba7e22cb8e3ca62a0dc1797aeb121e2289bbd7623ceaa33948e;
endpackage
package dat_110;
integer pat_num = 110;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7fa425768a70bf60cdc2e1488f8599f1ac32cfaace7103dc8636023a35fe38b56dfa8ea4e6010493142b2b0c5fd5247396479d1cb730e630275a423b231040a56b2f18c2a369459fc65f12ba31a3ca7777bfe1edb9e43106997de9fbd1e8f332;
reg [511:0] golden_data = 512'h78688c427bcce97475a54286ea2883a80d440e8be788c117f7b5bb4f4e81dfb4357924aa8cd146f30cb67466a4ca4e94b6c0f0ac1e34ec0ef642abfba149ac1c;
endpackage
package dat_111;
integer pat_num = 111;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7f995a6e4283724d72e6c2bd63df5ef580ba13bdbb6cc37bcac7ad76e5d297c376aeb032287346568195c33a49a5fd188e92840fe54d21e743876dc2a8f9c73202fd6200af05897cceb9062b5c7dc6155422d608ee1b17b4eed2576c98fd19c6;
reg [511:0] golden_data = 512'h2f2d618fe7ae6f08af032fd3b878dfdebd6d37cbcc2c02b65a060c796a3d042a3edf0eefe4ecb539ef65c71315b5607cc2332c7511888591cf4600a2c767b392;
endpackage
package dat_112;
integer pat_num = 112;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5bfbc1f8ccc5a345c73681856c704eb3487affbf8d88b7dad794391a9352517006cffabb056458b6fcf57bd55c880db85648c6dbf216be80cf8c831832debeb919306b16c21581bab7996c315a90c7b12f32658e24132ea50b7e4411bde88aeb;
reg [511:0] golden_data = 512'h666b6637071506ab2eec839b7c0079b9cf5a366d74f70d06fbf0c9cc3032559e485d29081a1b004ecfcad1ba16f0de0742dbe9e5e362313f437208c7793cfd66;
endpackage
package dat_113;
integer pat_num = 113;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h18ff6a4b78b55501301871afc6cf3f6378946f9f60ac171f42808763acb3ba5a041317fc6a4bcebceff7ee7b87d6ef1e8552f980d9a6ca18d53d77aaec7b28374e90842122c306f6e89080c49c43431e98870e4a4bd09d51563803ef7eb2733b;
reg [511:0] golden_data = 512'h6332bc0c98c87c7aeef4534d40916d11dc7151f5468dac1b1871e9c5c855c0d85194f1fda63c0f83d6b550c1575bb1679cb805b42723bbae27a9d61cc4d6d44a;
endpackage
package dat_114;
integer pat_num = 114;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h20f6b580dec59fed246617a0f94457e61d837b31ed297d83f32bc1430af174e02df1f127e537ea1498eff013f621b600fa0e9f703b1825a5e4d73cb45b818f160decd07c551e13a954b796a548961834fd8389477f5132f006122b3eb72199ef;
reg [511:0] golden_data = 512'h5f747c9dd14e48af70fc88d413631ff2a38daef1748d2bfb37bd9c5ec4bdb0a85c90f6da9b65b1b55dd11fdf50920a6adcf5a8c805881442d27601f2899c2560;
endpackage
package dat_115;
integer pat_num = 115;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h10b9da7c8fdec3f7c632821e699159e2c18ddaeb1d7253da1c5bd2503c484fa622e6616bc60edbd20b872fd3089759cd5680faea877fe442262a2d25b4ff0f406d7e9487075036dcd22cb3b6c1a79f6dea9e8cecca38d66a43546ef8fcc4fc61;
reg [511:0] golden_data = 512'h18e9ab924eee5cbfd330c96873cc7c128411fd9b17549dcb60e430295599ff467cd638a81e309c6690c7ed6cc4a58e3a4d98bd4fc7f4bedfa5243eae6ec7363c;
endpackage
package dat_116;
integer pat_num = 116;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3abdef3b5a7396964064b89533c1b9029bb389c3604ec01ed0aff3dde56bcb7d6d8eecbc4000713548ada379819b2175a3edffc4aac520c8a683e15785bbf9043ef2ffa200e5ae9cacf73449e66a6fe892be249687895429f758c92973a0e66a;
reg [511:0] golden_data = 512'h2730b54dec932b979586b7dd053485dddddf73e536720d7a79d44a035f51c64875ff6e6ae32e18626ad7f54a02bff3355f9bfa9244dd1397b6e7f2ac4ec55054;
endpackage
package dat_117;
integer pat_num = 117;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h52b4675b7360cf56183a3737667b71bf3fc7a502fae52097b557f916d889cf8b50e6428f14d8b4edbf5813ab4d1043e465b6c7a2f66a134df01dac26eb3ba07873b7a1ac02b6f429eb92a0b003011d1de67e1bf52f7a2d941e99f78bbd923f9a;
reg [511:0] golden_data = 512'h76a1fd26abd9708d3541b704b2feca65fb8f773592c2a1e88c1c7dd4eeb43be81cef9f8ce2c28a8e5d739cb9a4e1377ef097dec2360410323a69a582058b5dee;
endpackage
package dat_118;
integer pat_num = 118;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7277f8a60dd5d183ced83dc5715cd1f59781780c275fe093bea369b030a53df96d9bc2bee166ae547d7c2201cbbc6a71e8249775263652b86f63ccf71f809d084a59271b7c9272d4c731f634b9ae7b76a308f51e7f0bb68811f668cc62df86bc;
reg [511:0] golden_data = 512'h15163fec5c5d93b6c5b0cd90c2192fb99c4ebfac55665f81eaab379cc4563d764496583d582fd72b39ab5950e6b82cf288da51f8ab1a38ed7573ee2d60ef0f54;
endpackage
package dat_119;
integer pat_num = 119;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h37961499f0342797375b6649b122c1ab9df2434d7ed9545a81d0fd2efb9f8c773771bb16bd5c633c2765e4f3e52141060834879b4e7177e34cf68bf654f6f36556930e1e517f5722252a4b55869745f981923ce6d95fbba33a1cc4960405748d;
reg [511:0] golden_data = 512'h2151686b9e9708277fc697b49ffdf4c2ba7f3be6bcbfcf0852745e60d0067fee48ccab2cc7cd36a4db0ea8c5f0610fdc5cc96ac94214eea8d4c6a0dddadf9806;
endpackage
package dat_120;
integer pat_num = 120;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h784eb880e847e55bbabd37246f13a742cc2ce1a0ee8ff2f2af1a5ff6310fb2c31450ea0258b3c362f223efd984be6441e261c1fc4958552a5384cf91381209050a79345841ceebb8dbce3e2f030fb45eb6e2f2bfdd8658e4314a758c9810d1c8;
reg [511:0] golden_data = 512'h60355971d18c0adcbb5e59e4ccea06a7900a6acfc532de6786a22033407221d032e75b69cf15d61c9e88db67e4a46e4f4140d81c1542f1c07b090ab9151e9a18;
endpackage
package dat_121;
integer pat_num = 121;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4a6fe9bb458c9dc4321e8a091c3f8d9185848ac64a91c01fb19e5f051ab215d90dd5a8ff11523a9920cf5088212ffb9df8723b281f35590a9bd303e4d670503463f9d2c8cdb53e53c1b726f676eb65770f035dc0245d7a276e71545037bde877;
reg [511:0] golden_data = 512'h14624865203148d377d00a416848fd17af419f6a9d782271cfe3bcc98ab8e46c24e6f10d7735f84e38b4b050b34185535f8ddc8cfec93f68b36d21ce21ecd162;
endpackage
package dat_122;
integer pat_num = 122;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h59a8b4bbaf4d94c86dd9f84e508d06137c9a49c156880989749e688990ad381635749e2eba059c732130953ff8f8f40387c220882d6bb1f2cce725014b2c27d07a940a027021759650784a726a58e4fb197b8f8dc34c41b64cb5d32cc88fc4db;
reg [511:0] golden_data = 512'h1f654f314c3a7b502fcbf2e5e51a4c7890c11da5568794c4931052c9a24e0c6843784feeadbcc51afb933e49c2b8cd4cfe7a8f150250b254cedbefa393b1f0f6;
endpackage
package dat_123;
integer pat_num = 123;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7ea1c5a9c8c9be19eacce87e4dc3c0f311fc172e3e4209074c5405fa10c26426388c14ff61a842e9391a2aa698e14213721c880ac46b2c64d518e3b17f27836023e244a810fda1592c9ef385c5436d823004b13bda3717e26013ca78195a185c;
reg [511:0] golden_data = 512'h128dc76df7a7b5717185b54af9336586e1e7407f966feea247ddbae5d6da7eda6612bf1860869ff8973975f54a8c75cfa615754d123738255d9e5e926dca7606;
endpackage
package dat_124;
integer pat_num = 124;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0a2760a566ffc1948dc66b8357682176aa25e3604e3622fd4948ff92109338924351e078d52acc2d0a45de2abbbb43befc1f19b204d54f6a8b0324b5d67f61fd3b33c01b3b7ba5da73869ca901a34da97031379cdb7dfed59db8442ecdcd171c;
reg [511:0] golden_data = 512'h31e4cc827acfe89999214f237496a89b77ebebf4162dfefd2b7d85e74bf611aa41c1b73517c59019c4dd865e19140da0a8da01ef0e687d9319ba5fdca3117924;
endpackage
package dat_125;
integer pat_num = 125;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6204614b42b4ca73a26b9485f65bc5ba304278a2a57554ec6c1c206893ae3c14383c3133a21bebb77e7fcad8a3ab692742cf27656062097023c9ecf500971f5c58fd3bfb604f3883fe16b780476cdad6a771428bcb4e9eec8f78ea61bba42dce;
reg [511:0] golden_data = 512'h3f9c7e6aa1fe36feea15a0d2db44d7b31946dd26d2b528c130ff2c0d0bc4e572277c398e0ebec24a27b19b652e1ce4ab0c994af48c62a4b175bdf83d392d8f22;
endpackage
package dat_126;
integer pat_num = 126;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h63f8fa6c0364eb72bb45f5d9a201c85b6bd385ac231c069d2f489ce134f53da045991c78ba41e827d35ab7a59eac79b478522ad4e312984fda8b644e4b38c84d1fd44dee6d3e08b9475fd9c4b5a83abbcb3a0055173f13f1452f379567bfc5a7;
reg [511:0] golden_data = 512'h6e0282c2668d91773a90c78a8b64c08038f4162dc7e88770c4437ed99fd1cc941454303cf822590396700e59b56698a2e7ad739fa908ffe828d477ee12479cbc;
endpackage
package dat_127;
integer pat_num = 127;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h064479eeb253b8a1d813c135c4966d2ff20b5e342895ed0c61cc2d1cfccb113a7789e92b8a8465fb785d815ffcd66dabdcd3d8f312df22af16d059127e3ab2f0289c93cac207e643c6667e1a4c3113115a8823bbdcf191e9bb70b6674fbae665;
reg [511:0] golden_data = 512'h1d3b5bbfb273b85d0e2713ce33060ef95fb64050378128eb3e6605cc6dc9063a0e52f7dee6b74789cc38dd630f7dde19bf54efa333d6c54c1c76f6ce022c4970;
endpackage
package dat_128;
integer pat_num = 128;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h23d4ad4a907897128956424dc5330c23ad35a533005be4be0ef8fbc14d44078851095fb67eaa7b2383e4fb5e0543551ec811130d8838a07a8e84b02451c8acf22333d31a972bbd4378411217d5bad00cabf815f7356bca2a4d97f3245ed75673;
reg [511:0] golden_data = 512'h04c8ae5b245081d8cf5dcb647536bccbb02c40fc195f061f3b13247c6c04cf941b5240af1a95a6be3c8b5ca3ffb60f138586ba48578e562cd99928d2b65eadec;
endpackage
package dat_129;
integer pat_num = 129;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h149fe981312c32ffff798d73862fa7c2b948e5a4ff27594da51cffe9dee933c62b445a84843a83ecaef32e6b9387ec693599fb2bef33db236dca5358ecc2e5511f425a56edabb1ab86adfaad51b935a07f1d8c97a070fa57ddfa22969d34bf97;
reg [511:0] golden_data = 512'h66063946532146c654c126e01989acc9272be60a96de74bf010b3324cd85c544646c018abaef2c2f7555cde782dc21a24f43e68b3474bf57fa5c11c71951e484;
endpackage
package dat_130;
integer pat_num = 130;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h37acb0078b1e1d63a33821eacc2553550d105e30d3a44ab4e909f31e690ff66c09b179a946acc0cbcf350816f60fa4b1c4a744496d9eecabdd155b80bdad5071104a5357037aa23cbe9382a46f5a7422cc166703b5e4bee10c6250a1f53bd65e;
reg [511:0] golden_data = 512'h7fe086aa127472a2c7b459b7e825126f82cf2f0464c0a109e8e3b7cb4a063372561270bcdef2933f8b797a15dffee610f398d53942f695f684c8a3b620d39088;
endpackage
package dat_131;
integer pat_num = 131;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3891f0a01a8e8dbbd0cfd6fe3808b5dfc058abf05af86e5dcbc9fa7166898afb5eeb841149c825e751b356655cfe516a1d588f8e16a837aa3511af68046890a31d11f725fa1e7fce5cd5143fbeea478ba4031fcb08e2524f1d41d4dc5d645cde;
reg [511:0] golden_data = 512'h6b873f5f6397a4a31435d2deb934d82ad617be7c1637f824447ff7b299c1c64a68e531a0e09ead00513b3850a342d238733a013bff3b8c47d0a1d471aaccd0be;
endpackage
package dat_132;
integer pat_num = 132;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7540781c53a72af6d1b986436254844c98b97d00edb3d1cf3a3cc5513f7fc7767ca45d5d51996e4b0e2901f59eb7ae780418161af973f958075160528d442d0044f55bf1a76f7a6dfde8fcd85e1f3a6d5cfc0380ebcc1c229eecf6a6fa20ecfd;
reg [511:0] golden_data = 512'h5a16069208be8889d938de46b3a439a86b7d94ed2217edde48ddc0f7642e5ada1ea56f95477e5ba8a33b170e0a20f00d21ebf90e4218240387fb30b19a5b1a64;
endpackage
package dat_133;
integer pat_num = 133;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3eaa95b8bef69ef34e4e94de7281cfd10c0f598cba0deea5f52d4618c867445d62830e0b8a4315d199445a4ffda99e2b780225cc6ef98715484ea1a4e9ff633016a088d2798bbf5c8c15c0ab24a495c4d47b2de00ddee6e2de21141fc76811ea;
reg [511:0] golden_data = 512'h0ce4add9eee3d10855bf6e1db019866adae67ca2342043b9d45d5aaff5afa0b04880e253252c26c0a6893be38f59ebfbd46345a2aa58241cf3832ef2a4764698;
endpackage
package dat_134;
integer pat_num = 134;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5d51b9ba0487ea9b73022210b7d654a8e106d7f66d06a9898184e6654cec77784c70a43ef366c36cb699a104a33bb7062b26baee2585e36105855b3286fd83f047318ffea54b16fffa2e38b80abbd3e113a685796d53afc89bf963c776c2d22e;
reg [511:0] golden_data = 512'h4a7291231a716b99afcf676474e259245ca5579e97b877a4bc1a80167e4f426418a1d6925d36bda55968abee1586793b25db4a22368fc5412d9841330ffa47f4;
endpackage
package dat_135;
integer pat_num = 135;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1d214b3740a6aa996985b72b7235840510143694c95a26569746e0de6aade5d70cd5de45de82201ec038cec55bfcf461c4a9858a724005a6a90e314a73e650c059dcad452ad2c809a9d210d50393fbd9966df961290f2fcc1abbacc5ff1ed120;
reg [511:0] golden_data = 512'h5be0996de1312be49955985e610bfe955d5b49a14136be8e8877b60431f3cb521d8cba9e93ea088b0ae470ffaf10ecb0804ba8d0b1f64d7d7ca5fd5fb52d4434;
endpackage
package dat_136;
integer pat_num = 136;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h50755b0c6bebda199dc1304889b9d43748ff6adf21a84344353a63899e24d91d720a9ca79578bd76b91b3df9c4f2021089e7c2179ddd294d891159b7c94392627e08c74766c3a7e0cbc0645d60935b1344bfd8fd69c83d5e714e42d79d232b59;
reg [511:0] golden_data = 512'h777383bfd0ef73b028e4a24af8cc92467a2de022979b798b23749ace614dcc9c2cff0acd0ed810857a15c220d04e920e58a6fddf45b59b8f2d29bebad7c27b72;
endpackage
package dat_137;
integer pat_num = 137;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h04fbd9a136946cbdeb4dda0e660317f8b0fee2c23169c00f9bc18c6ab25671ac7eb831a9907d59543dbcbc7aa72476b3150c0e683e3d0062b08cee7ba1d4cd3c23d9fe04c7874c19c59ebfd3216474add6e3ce6cd334bae939093997912ff965;
reg [511:0] golden_data = 512'h446b5f81dce9231b9cf782354497531c78fd60cfaecb7f68e149edd4f4fd70a0611fdbc74d62d99a2a8775089e43dfa587c05d847775f7217cd892e9831f5bb4;
endpackage
package dat_138;
integer pat_num = 138;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h512be1ca593be27b2390e778efbb0257cd6e9c989b8ddb5910e466951e24061e4e8ae845d7a95d2fbb71c8fec80e70efbf4e7c627a7b5fce705db4d9d491d4701b969d48ca8d2bfc435a096886fe2ad0072cd212cc3431104ef2f2593b3e0998;
reg [511:0] golden_data = 512'h499daae040ac685c1cebe0490d964998661087c42812a40b166298d5807e7d7807da62d903652540eb15a64b28385a8363e16fda3e4e3d035148731b4578eabe;
endpackage
package dat_139;
integer pat_num = 139;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1b7fd0df39424cca4a950bff583ea7ada4288164350e08722ef84f80cb96121b3b3689ad3b9779ee6ec6c6ffcd64f96e10829d5e585c09b641758dd95bea454e76555245e9977491c8f37859dd407a70cdaa146df0dbbf2f45531bd30fa6d4c4;
reg [511:0] golden_data = 512'h1e5f48567dbcbf6d3db28cde149ae4d0d211118cc1c6189ecf405a81215b94a81f5dc003fa49674d854cab82c7e549a6c899a8bf24bf4e91b7f9eb47e46ea230;
endpackage
package dat_140;
integer pat_num = 140;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3b2ff4430b11c05538a0719c94d1f0a2f0fa08afdae75f89733a605889c793756726544e5450c4715d2dc0661e503e499ee60ac824d4bba090a42a3e0cc04b5668a1973eb8ec8e4fa6ddeb33c1d5597dcbad9205ca9c2f7a3bbc690af457cb5d;
reg [511:0] golden_data = 512'h4a7ba191f6919771278fb7395ca9085acb03406307b5ad4831a701160f2eb53a3a2f0fe8553f105028d22d8acbf9ba88f62faff848cd614a4982020b33c7e57c;
endpackage
package dat_141;
integer pat_num = 141;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5f8e96ec5ba3582b3282071989527e211a9036f9e32aa1dc893f3fc12830700d49be303bf9515b328d9b351ec9e9ae7e131383d918246dcb55b810d9c3e4e2df36ee2eb22a43b681968bf6ac792141425e980dc9ff58d0f986193303da932dcf;
reg [511:0] golden_data = 512'h2c240cba24684a3b13a2dadcc9bca63013c649b37784111f03e675d9fa7feb960bfaec48b766ff825a94be82141d97b08c7752ab144f60438cf55a3f918c8f8e;
endpackage
package dat_142;
integer pat_num = 142;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h689925adaca75a6175c02a88a1421cdb7e5da592c1b2f41fa846c39a0e0eddce20fd4c2a63b1176ab8f664cfb5764fde3c0f41a9e3ba1f008e017dac6026a74d68c8b858963a9b2696a87554097781ea0ad81393d646c3017bfe74cf13683e4e;
reg [511:0] golden_data = 512'h64d0c448f8dd608c7eb1bac7e2c53bf9d5ba91b08754cb06b1e05a164a34501861df9b6fdfe0dce069b910510ac385bb8d28ace1bb7497cc58173f7c7f88f7c8;
endpackage
package dat_143;
integer pat_num = 143;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2ffe71a3734724ad1159d8ad57f0c99d0dcbfb4a05e989adbd1a043af9f494e80b796f9de9d4bda7985c01b07bdf86e4012f51c70953fd7874d48050d993b0717a80ff68a849a8318fea09ec5abb846e7ee54646d5d7143c1d115010649373d5;
reg [511:0] golden_data = 512'h7ff9ff1cf5ebabdcf3f9a4e32ece253a8ce04dd0b0796d8d903b8033a86a741a5a2124fbeeb289ff61056b9711490edd6e017e9d52c23a764fe98054639d8922;
endpackage
package dat_144;
integer pat_num = 144;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2a834354624610af3cb017a31abf47f47bde710bef3ea2f2475edf15f58ed42c3c2374423842eb8fa26b5b14687e3a05860ebbcca5077d2c627c09ae79db1a8761e928e31327095c25331aec6462818ae678a77d4da0f67fa7fd408dbd5945e2;
reg [511:0] golden_data = 512'h0ecdba9669934cb73b936c7ecedd93880911d7f7531d6463668e0e091d29b82874c1e914fde6e269f51dc92d49a87db513fe6c3c21f6a2f3eb00ed11ea3fbe86;
endpackage
package dat_145;
integer pat_num = 145;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h325b3264c5d77ad5a6369a1e2f25831005177c45429374f595e0e203399ff4bc0af0cb7f1a7000f2928ac8f01c036d98f418ecd3914efa5a5d7c514da868fcf03882ae8e07262680ec868b660b8155420573bcdc38d897729a75601efe63b036;
reg [511:0] golden_data = 512'h556cebcf34b52b069bed9ba55a52d904f3c7ef7fe62529d9a96a02c068692dae64fd773b79f1705311c92c5b7c6b7a307cb5b427c4b32d03c10966f6d08c38d8;
endpackage
package dat_146;
integer pat_num = 146;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h280f15d94703d3d0f0da1ed6b6b9de6e5cd1eb28067d02b75808ba78d7e461c01e375bbbaf372c348bd79c7470e2ae8ea4b81ad46992f00599612804288af55c08e7501b912d6f9f510c081a9632772c44f759a4a12677d5c58f9903715476c8;
reg [511:0] golden_data = 512'h4e1e39e14520720346ddc99d9a0fa5b751ebff60c8550fb39a89a08c59377cf87f51c0f0e0b5c0aeb77ca8a3120b92d94f9fef23bb2c0fa78798930b08d0d058;
endpackage
package dat_147;
integer pat_num = 147;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7feaf305a9eef891851bd76f226ce44f393ef62f8ce5aade1e97fe0638f8c95e7f4ec199619d582c8cbae5ecbc9cf07adba754c76d040ddacc28abb09b4b674101cce493842ef9e1c18ec69ab2443feb765a132c94d71ccd92e3268471f5a277;
reg [511:0] golden_data = 512'h11e97bd959f870372cfea63cff5041dea5c8463c9b85caf133475e46be2222b07bc716c1b1dc4a535e22b85263dc60cd410e503e64c3aa9f603e7fc753942522;
endpackage
package dat_148;
integer pat_num = 148;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0ceb7d13d495e0436e72e13039a2fdf7fed81652371e8e1f84699601f1f333550fb01904f312b911547c7155a95cd0f73d31eb125e8ae1ac7d069f53b35418131fe857950c100f6ca075549b1a4387bc2778888ee9c143aaba39ec0773134fcb;
reg [511:0] golden_data = 512'h6471a21e428b3d1ba58a95e91ff04d665e1ebb4bcd894205942f5d671a51149232b65799c955482f6d438f9b9d043501a47366c259f71593a32ca8087c9a70d0;
endpackage
package dat_149;
integer pat_num = 149;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5f562a1bcf3d538f117269a3ddc4e00dd2105b3e9a5f433db0cf895ea0f36da309d9d3aef74081e1522d0bfa0a34c74ee5ff49658da68d3d17aadbe6a1f46922576816930dd32a52ecc7e8e9b8347851de3f907830ba1496f6bc63b6283d1a59;
reg [511:0] golden_data = 512'h44842835005bd753ca38e6ae2102ad4aa654d673cd189868e6adabdffc6d8f7c47e94f20335c4aaebb84e83edc824e128a7f42d537c8fd9f7a40fe3d7733f12c;
endpackage
package dat_150;
integer pat_num = 150;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h00d65deed89d50629a827bbf94c96ae0609e79fc81981725d8db3379421bdc47141b00caf12438ac652261365aaf35cd7a2e6310df6c6cb154d787bb9b9f5f781d91a04df74c71185853a2e7d29f56d0c55b3cc999170c514971aaf7f85a919e;
reg [511:0] golden_data = 512'h7e3c093b0efd6dc9491e48e23be9bfaeaa9ac840465e80e7b37c481210bb36b279f4ada327b4cc2d4f35c88418c2fc8e0f8776128c55e331ed4dc62a3308e38a;
endpackage
package dat_151;
integer pat_num = 151;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h038292d212d650d8973ede65e7bf5af77b44a7c2b8e3376b803a896df34b5b4a3829a508d72f9a6debeb7ac0bfe99cd6e334591ccd0ca7b4cf9dba709d2a398b36052d45f65901da629fc639889ac04201b3a09b31957c6604ba0ebf9cd7871d;
reg [511:0] golden_data = 512'h492e8157efca40c72cda636a6cedc9c2df2f6289a8b0abfb9b30ec63ab0a442a2a780000825601a722459d5950f024507ab0b2e8e83ebba5ae4e4474fb6df5d2;
endpackage
package dat_152;
integer pat_num = 152;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h16956d3883942984f5c6c6d987113740be62fa9d73c9331eea90be7392d1e72b45795cc39d94b770dd8c77ef5ceec20782a3543ef756fda8f2f455d07fa9109d7970f4d16b184889508b303e7ed2efa9fa392a0296bd3bc35cdaa590ba1315c2;
reg [511:0] golden_data = 512'h5923fff8f064010c626bc16e8a8e3db558d820278768b9f8430a1344835ab518617b2c0068af010d1fa70398c6d464855722c02b25639fd2a24d109df8baad16;
endpackage
package dat_153;
integer pat_num = 153;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4dacd0482f063382a491409a04ffaf6deccd5155eeab291345e3f952a381c07a0f62ff94e14545849d237943dfca0db837da5890789b0274f54efeb1b0b43afb7dd38d868103136fb9dcf84287a2ee17e46b24576b670711ba814a39ba988145;
reg [511:0] golden_data = 512'h68f0bee5de1a2a12bf4b233c38c929083e254c55c5920228c237cfa452aef0e20fdd20a95fb6b8c6223ea58be7db033775de68630eb6444eb17bb3942d10147e;
endpackage
package dat_154;
integer pat_num = 154;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h616117cd3713465835fd147bc39fe13bc6c092e5122a59143e4d04055fe158610d73e0bb660cc2e7ed7a0b42366094c45ac0f6a52b4c360912456cee3c10dd54324c9f6b0631b8b39d6485a078ced6638ab3d945bb5219c9b02794f1422af0f4;
reg [511:0] golden_data = 512'h3fdd38bac62c74d409a33f23af439d613d0d278e24fb6bcc71b887c419cb2ca0213a43bc210fd582547f4f7da50f498966dd8e924421907dd73f79edf4836f5c;
endpackage
package dat_155;
integer pat_num = 155;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h72eab1dc10a1c3f9467d76d332bd72ca30f511db60116c525c83cbff21e511cb3b98096e6023dcbb5f61c9eee7e34a33bd57dd54b7ec0f62543458e35787f06377dcd9feb05289e7651ae03af68aac0b01c58c698db47f5e427ae457b5ec76b5;
reg [511:0] golden_data = 512'h63f100c5003a20cd3f8b7a6a686ffcda2076699cba266a738b52169a89e73cf43ec023d5ab493897ce82919708c8644fc6a54759c1a2e15704bd856545e511a8;
endpackage
package dat_156;
integer pat_num = 156;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6c9b5646c0941a6a2573b932d814c79535e0cc60c83fee9942ecd5377630f4f04a3cf084b8452f12300308b11a23fb52be8a7bb919f8b296b3b0628553834d6e2a148af45b553c199ca0c8bb61e29ff8fca5194928793983097536fe03be72b6;
reg [511:0] golden_data = 512'h7fc11da5cdd6931c7754a15dd03d05c2ecf8e76578e26c36d1d988172fb28afe74a4f41df4a533a7a99e721ee7907e77500cef1301931397870e4d15624fbcd2;
endpackage
package dat_157;
integer pat_num = 157;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6ced37127824874f17eceea0dcf33a4ad1371b92a823672409951182d58e031576ed81fdbf7824af284c47a77143d76e3b83ec1f9924d91b46959c98b662eae07abf2389efcf1c287b77e286f74dc66a8d6ecb88e444b3d8f7b4f93910edc16e;
reg [511:0] golden_data = 512'h58a04a37cee37dccf399b0886aab69c37aeb118ee602a79e5c1b80b53f2155665c724187dd0dd9fcd0527b637e400851bc92f91d96c7edbe2948523ca8f7f248;
endpackage
package dat_158;
integer pat_num = 158;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h18abc9d006704c506b33eed564bb6d3c35ca8eb86d2f3b4e59e7fffcc75334d61dac92bc46c463532d6f8780e6af95ed867748935b51e0eec30a56a3278a9e23453ca435dcbe3270f864512f50f3c68f4bde9835cd1490f381fa88b3570a436e;
reg [511:0] golden_data = 512'h13298f5c1128d907ab892a2159b9c1a3fe3aaf203922f6b1551e731ffcfae1a8578c307f7fdbf332c79cfce61ee3faabf478b0692b3133e8c07f745915335d78;
endpackage
package dat_159;
integer pat_num = 159;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h352c840e9cb8cadafa53c70f0989fb1dbe14b595d0761a0c01a1f50dc0c03faa1426ac1d7dcc016d4d1f36248ac2dd9984c4d3138cfdf7cf2baefaf664cce9c16d6f717bccdf12f6877e164808488c7bd8a52a9ceefa5097d21ccd159f1f64b1;
reg [511:0] golden_data = 512'h2d46030bc699b84be7d89fa2654413a1dd0b662a1eb836cb22cb34704111284c5d5db70e24ba54e131e4500e08a62ea05f870feaa444e62090abe7ab008fd9d0;
endpackage
package dat_160;
integer pat_num = 160;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h46c30dc073fa19652fcba9a65171d210e9f924d9e693918faa9b3caed9e2682067bfe1c11d5344cc25a64167d35a6fb06a46a42b59d7f41164294da952eb2faf30447f5622ec94f0366bd09f9e86cc62c96efbbc47280a02c4c9114b81413ffd;
reg [511:0] golden_data = 512'h212a19a141099a6467c910af45351cd2b31925ead0c64feec39406561058f3c67bfe7f72b5347463890b69aa79f06de0dfd207098d2d2df35c844ae7408b70c4;
endpackage
package dat_161;
integer pat_num = 161;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0a6c67405c75b5bd80e9716862063f3a5aec48f9257d9cd120ba49a9afd269bf502e7b4a71b8a99d3e31471c11eda0137ea9d2fcbcc8ee641c14597afa3439b76ee5144c0694fdc2ef597f7f8b2763a14e2f6b9c72c15f842a547e4edcdda27a;
reg [511:0] golden_data = 512'h2ce4bd31067420b4eedf456a2ed02112528ff3897c71f9d38198fef2e924de7a69e30b5cd1ab8b3d5ed31be2c0894a7d9c8ec5c5703086c7fcad4df85ab0e26c;
endpackage
package dat_162;
integer pat_num = 162;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h67e35db422c508395fee7e9108ea0d390cb7213fbf8d8cbe718d99f84311646b4efcbe8300335b311e611529c6dfaf87df80308bbe8d95fc77f7beeb34fc7de85a8693340a694e2708929fe2ea05130a20a8ea4540bbca6e5af37ba92785ecc3;
reg [511:0] golden_data = 512'h780769387ca045c0a6ac55db11cea0882881057bc0d68c707bf3e7c556a7ff704c6255d64af80a9308194f9797052835f03bff3177593d6b115acd9cd6605982;
endpackage
package dat_163;
integer pat_num = 163;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h24db7b137ac52319575b7b449d42408c5183f5afc6508b1012647ecabf96a68d45db2faace5eda33efd6165aaf1e79b00bbbd14c181b257b762b9a6cd33ce3e61cdef77c04a27d7d3aebba6ff8c6618f48cf04ea42520cd7a8c870abfb88f2b3;
reg [511:0] golden_data = 512'h557956c7f850456e128bdd4e6e79203052ba4116106ec884acdc0112e469aabe64c595a58346f97aa35a3b56cd288e310c852ae09e5c416c0168852afdb4db96;
endpackage
package dat_164;
integer pat_num = 164;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h47ac811a9b91aabd1f1dcea6e295b3d99df37023f36210f4784e2ead0f7312ad4c5f13f6366642e91f3e40b01d1cd7cc57e549f28b6011b623c4c9188d1f449307fdde785f0dc6f255ef449e6ab1529b16ccffeaf5b4af59e117bce0dc8a56d7;
reg [511:0] golden_data = 512'h01d58b3ca18a6e7601bb2426cb9bb53fa4eb7213b71576ecddd8236326d6018479daae6a99973f0223ac417f66c007ff905cb87e6e753ebbba0ad3e4548ac636;
endpackage
package dat_165;
integer pat_num = 165;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4096c6fecd61df721c9cf4706cc4456865b17a8420d3db36aa34ee92d3d58279357a762b9385487718dd72bfa45a63edc8d728f5268411c6f8edb287b6aa860f6ec7cdc7c5ee12d886eb296ac13236f07ab112beb4ea6c860492e588f9a3639f;
reg [511:0] golden_data = 512'h702ff47c655149c8cd962bb6f9baed28872d70ae305b1a40ef7c3d2a88cbcb320004447224bb46e71041a514a6b540a793c324a812d8d8dff4315b6f308db4e2;
endpackage
package dat_166;
integer pat_num = 166;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h50bfdf57fce8c0fcba44d4a0b9775e2cb7d67f9a4bc4e91ecb6972020331760d049696b6b188935b1dac016b661e70f1c7866f9c57af676b07623b71d138f4697ca88d4a9d80610952151c8e12d5798227a2b44721e6b5abd72373d6dab5405e;
reg [511:0] golden_data = 512'h0b23fa535643d43ebb47ce739a3ef188e2233fceb26cbeeff6588429b44bccbe54204b8085d3279a982fdec754396bb2b121910b645c47031c1657edfa435dca;
endpackage
package dat_167;
integer pat_num = 167;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2b5283fed9c0a11e0ff29daddf4adb4c8e4427d256af173103b282d1eb207a765657be457cd2f3889aa61daa9597bbdaf7a6df16f184e9bfad9e4a55a2b58b4e792a95477cdc966d82180c7a8b801efdd672bbafc7105132c0c0f107194c7a0c;
reg [511:0] golden_data = 512'h0dd856fdebda2ffa87456e3e5f7ed23778e1c44e8321e97829ea81c5cdc776aa4ab2b78059ed53ee2d9aad2938bfa032c400c7b2f6906f9d9372b7015a17f7c4;
endpackage
package dat_168;
integer pat_num = 168;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h64d5c2c22d936d75009d5bd8bc65bcb86e7db30c5faa21e9857b436f6e4eb05334086cdea133d80440cc21abb772b97c4992cb207cc1d60ebe0aa33f2dab456c3e2d5f29bd07df0de4e4794e7c0cae4d38136d968ab7dff31e4acc3b7a0bd671;
reg [511:0] golden_data = 512'h7711b80659288218ddd13ff013ddd976c25d82de848d52504a7fd76fe02ab6aa1105d65b92805d9eb97fbe55944939fd2a7d08d2c3ee38620b900b832a4dcc20;
endpackage
package dat_169;
integer pat_num = 169;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h40122ce6df54c3381afff06213955f6969b0dd97bfff8dc8065b2ab30992dd0229593e2a978165f2e345d3b3176b5d7987c1d7914c3a548fa8ce5c8f9f8902226f3df172afd62dfa1055dbb84c7b56182c3f00ab8c9523cd29217d4aa79fe38a;
reg [511:0] golden_data = 512'h1aa01696ddc6232e4e7530f5d3d67b592b245b67719a048de980c203d6d4653e3e1c2f519fb4bd4e35a60d6009e780b746e7e47a40ba8cbed5188f93c13107ea;
endpackage
package dat_170;
integer pat_num = 170;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5526017255e95773cbdd198e96bf916e7687c9d9087c05c7524e4d0f9bc5c325171a0a6210e767cd70ea9684dca69fd21fec7da0c43873b29a8708c8736b2a2730b5e5d09952a7481abafbcd902d05541d1f8c1823f01f5769b7fb4798158d73;
reg [511:0] golden_data = 512'h5ccab08a4d6098bd60ab696e70d5ccb89f4523ad053fcba54e5ea16af2380410327dbedef5709b07ecf93d68856e368fb4a92c13c415b01b1be560c624f31a1c;
endpackage
package dat_171;
integer pat_num = 171;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h71f12ea43bc3c28b4d76305a54922ba4d541227f6616287c51223e8a3a0a8e266b5deec2e5a3d940692e6abf3376dfd305a45960d92775678757ce8f63cba5d75a020251afbb66c61e5ba70de555d36d750702c1df1bf430cb0c74b89f3b6c97;
reg [511:0] golden_data = 512'h0bf0029ee76747191279decb909481c050a03f26135c351cf0ec4faf94056a8221e6ab308dc4926f58f0dc60837959e207038de38d8bd23ab7e9917c8ec78aa0;
endpackage
package dat_172;
integer pat_num = 172;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4e4c8626bb50f4d2eedde4bf36a6598fb8a091683a0adb863f50827681622b953ee72af5c1aede3a780bebe4772940c2f1c45ef40ace0fd2826bc73e49fad6b551b2d48c55de3069b3e0e005c8b292728ad477863ac75c04d9fcd1964d479252;
reg [511:0] golden_data = 512'h3f7bd9b09e38077f387e3cbee491e6ed11b1a50d2d121e332a1c827e00b0eb6667ee34d06c903769307eb2250b8df8c60da012bb2c187b85247d880351b1cd1c;
endpackage
package dat_173;
integer pat_num = 173;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h576dc020191656e16bf8f038a1da0179a57ce629b3aa3fcbb128524377756e4c1cba869e42f8f44acda2a72d0a2a7f6f1bb732ad2f39ff5d61dc33824b8f58ea5e7003d9ef4c0f8fba29da2486565ca62ffd4392967073c1c28c0d339dcf2726;
reg [511:0] golden_data = 512'h7580d8f517363e487447ec8dd9b4704307a4e09b6926aa1b6e226d7eb30e1a5c6a2c7f7ea212ff52d0e41610afbebb3792d0204c7b3fc6e68bd8682f7e71c7fa;
endpackage
package dat_174;
integer pat_num = 174;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h272df4a9c24091214c4f4aa4b9c63cbc485cce2c4b8daba286fd9dc14c937afd7992a4f1eb51d95e8ff823ee7df811c407575a8a21d9ebfea320ba0d2d874b9e57f143d738b98d22a7991122220994ba7974e06baec40c552fdf6f2dd2822142;
reg [511:0] golden_data = 512'h663dbd6373be249c8e5db69f553f781f2bab0cfcfa623186c92f3c66d5b2fc1e302c15582a48351f46e601748b152fb4967fe7b149ef4b8f10f5f6e523dd5b90;
endpackage
package dat_175;
integer pat_num = 175;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h18028f8348c23562a22552721c93e0d04c1cb9de8fff97c8d9db927e45bb6cac1a96e340f108441ab6dfe3930b6842bb09050e02c5deefb1f4f931aec9bfa3b1751f1c259640ab88732c0efac48be3fcbd4460b8a589acca3c32068d9df2c256;
reg [511:0] golden_data = 512'h02b8cd9a5238c28ffdc745aec71d4fac1e7618dbfcfbfc12356320519a5b785e6ba9d36a1f9ff9eb4d0e03754328d9e72f17cac52f0577bc4a0d191895f1e610;
endpackage
package dat_176;
integer pat_num = 176;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3835afb752efdc298a7bab0a047674c3b3d467f58ad283e3d888c38a06ca021161491d0c7e1b19a5110ed6f09723708ec027a2bfac8b818a25650994973830741c70f8fa973c37540177af61ddfed1bc55e061c429bec45824f4544636c0a4a7;
reg [511:0] golden_data = 512'h34298c5a2199ed375c0170b5773a753ad923c575d84f04394a29d663e55b9af443e049265070101cf48a0f4b61df6ed2c86df648efe7fff5aa38c38471ed6c8c;
endpackage
package dat_177;
integer pat_num = 177;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2972d12c37a99c1435e6a807952954ff9c27d90c6e2d923b02ceac6c5a20642c4ceb1f92a31274ef7d0ba2fe627bf45417da9f71592370be84c876639cd0702d12ea335e874a842a369fa367e31bdcf405786d1fc2b6a266cec6e3076201c767;
reg [511:0] golden_data = 512'h0fcd3ba364e8869f02705c836a523e3164146f8007f8a4b0c5ac6fe45e776f4832e59240f1b0648aed30268ee33893671bc27d418a8a8d850605a7c62a4734a6;
endpackage
package dat_178;
integer pat_num = 178;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2c390b64e0d59a03fe5513f45a2cdc179b8d13a8265d8157724a68a75a467d4c0ce62b558162e3e30c12bf5e6ace9afccb9cea8e6b08604d8f21164c9a889ba55306ba2b3a4c04f365ca4d874b6e68eb17590e47ccd420089863b6a2878471d2;
reg [511:0] golden_data = 512'h6eb3d597bed9d1c0cb4cbd6737fe2fd50d758e95568b2f5cc3945930f08c52d0337b6cf593fbed73652dd8a86195f9a710cb6b63cd338bdd454e931a763a65f0;
endpackage
package dat_179;
integer pat_num = 179;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0ebc01e656b5a0fea045863c7a4f8c4180ae6f050fe27463b2182c8a835a36ab2f21497c7933ac457c66abfa1fadfee9d308b7763d872d6e0db8baaa6e733ee734e11efcd4abec1301168fa69743d0ce01bff1adcbffa6a96ff1e01f59549d90;
reg [511:0] golden_data = 512'h7a69bd8d8afcbf718c892b2b7b28ae129c4f61edbd7b45dc6f872def439d0f741898634b5e51fd45c3953cba232f88ddbeb62758c649c240302188952ea57bee;
endpackage
package dat_180;
integer pat_num = 180;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h00b87544ec829b34f7e14a1f557202edb678eaf10a926d8922447893c17ef42c532ec5a36a1326e1161a019db9e74628e06c05f0f3e7a5ec57dccf71b713650b3299ff1f19b9356157c66273fdeda80c7f9c82a88f96836d89cdf8d755412d7f;
reg [511:0] golden_data = 512'h497b74c3a19b80522b1099def8bbeec31d67309428291e0336aba7576ec6252c76bef47983076ea09b6c727208adb1ab42511fe675eff8c166e451bb82fb68a0;
endpackage
package dat_181;
integer pat_num = 181;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1a9566662d0d85b5029b0f008817001cf9a16517c16abb5c2aad8e4e8fab5d2077bbc8a50962feef74dbf68a4ff74007eea8d61a75e3891c6707c2dfc3f8b7ce622749904890effe72346bccbd3f36ad0fac2e04c5467ee8ba081d6d036005a8;
reg [511:0] golden_data = 512'h2dbba9b1d7ff6dcfb0f33cefa2a3e59184e0a33c230f43e30c2745386248f95e55ad25d8f2acc89f0caf27e129b2298df8962dac61a59aaa24df259482192b62;
endpackage
package dat_182;
integer pat_num = 182;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2d22429017b47f9bf0ce5678f8498fb4644e57877c93485e388ddb24ee8eb62937f96416001a7af5ed0f1b52df573071e5907b3145bc0b973c152adfb522e8636603332af439fa3b81b0f68d59d0df2e3f842eb5e10b6f15db698b1161ac1567;
reg [511:0] golden_data = 512'h3273a6279ae38dc7c8d5036259ab7555d55438cd14a607cbe267ee053601240c32e066277a2efdcf04e10a1c04521ff94b4963079da8e05074ba7495f4eb14f8;
endpackage
package dat_183;
integer pat_num = 183;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h102fd382ba733f867bb3e8daceca02290a18c7813e6bbf9e386fffc95e3a26b45a6d56271bd107518f4d8161da9804c467f5a52ba9302315212dbf31986cd9c90d09f307e6d4578537164424a35d7c70fd3e64d040b1eaf2d5eaf6108fddb0cc;
reg [511:0] golden_data = 512'h6bce97dc65fefd0b816010019e7895b0d6accc733a7a139340244ae29b7722f615ecc2c7148d998ef7ca11d5948abe909bcaa16c5afd31e815446b8415c51388;
endpackage
package dat_184;
integer pat_num = 184;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4c476c3f91ef1a117e89ac9805bd6194fcf8795da5a0923284db8ca1d3ba30ba073b4811cefd0cb6ed30bb3a07e85c97ed9ab4a5d68fe9951b056836726fb43538e11060d30fa6dd82cf407c3af0d6c76b29b35652bd1cdeead373f8b1e3845d;
reg [511:0] golden_data = 512'h4605267324678861f3d5fa751992f52014d7874a124d469ab894716bc30017ac6348a40f07eaadfaa043eb60d054c064247970aa435d40d49a4eb038f54e2faa;
endpackage
package dat_185;
integer pat_num = 185;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7815b957c0dd17764e01c04e3211feffc025ffb9d145d6ef3802e1e5f698176a350086b74930a09bb9e878a5af45273d55db44458905a6da59d297f7917bae063b6d76b091385ea47a45b5d979183863e89260f7fb1b79c9134e09c39899cd45;
reg [511:0] golden_data = 512'h6a9ecd32797fa0d98998f7ebca6201c2d43d17a8a21c79697748a0c56f7091a269902eb9d0ed74b18ed7598444b1c9078f8bb04e25c9766de081828d170f664a;
endpackage
package dat_186;
integer pat_num = 186;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h770a5cb7a4f8a27145e1208b8ebcad3f1a29dc37f6428d5b6fa0111a0bdc16e51aa229f260bfa16fee5b8664c0fd5408621818e9c963814303490b2c89c40a4378a1e978e33de9afe6d8e9fe06185a3d2cede9bd6200423b62852ee939cac180;
reg [511:0] golden_data = 512'h2da812fac797b2a0fa99aa48763a1f3fb9514f00fe2193a1085772d712f09ee634b129b0080209ba3513d5a477d367b03e295e73ec2253e5f1a81c56336db9c0;
endpackage
package dat_187;
integer pat_num = 187;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h74f3528155aee6412e269fce908b4ab210d960641703d1b42d685fa14eb2a4823a9d9d336b0021f522a379af47fd8c9fd3299213444a8b51867069a5e29b29c04e96129dbd0c38ae4f035be7375ddc3867d06a64fa64b32ae9c9f1684ce77609;
reg [511:0] golden_data = 512'h6a4f0236db514becd30c2c03dfd68275fed9ef14b22662f4bcb23f6dffd6e2ee6a821b21d6cfe9120c6548a7b89446df827864f87032ccfe2df9ed588e10eb58;
endpackage
package dat_188;
integer pat_num = 188;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6540bbc1d257e66903da4cd629b270506d36e26ac72e2ba212ce3f7fdead1b9c448578d4990345e2f234fee3b4db71db453f2a6dfac955b348ccb77320c6aa8b4cdb1c9dce2598b782a8ca1bb0ad063dc0a2d261c0e14f94528107b31fe0bb65;
reg [511:0] golden_data = 512'h4b2aaf7136aed25ed4b333ef010b97077a2060f1f1445e517840200fe29e3aa476cc25f2e3941564c8ee68673f400d6454cb58b878cc59987ebb8fc69591223c;
endpackage
package dat_189;
integer pat_num = 189;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h65a11fb6bab9e962614b74f580fbf4fd911a50d084379b988feeadfc04e51d6c76fe57263b430915d0064db6d718694bc865f83c2ef5574a8965c6d66e70744f3765818257b54ec56c167cd6ee0a1acd8fcecef81dabeb595a6b7fbb92d27596;
reg [511:0] golden_data = 512'h7c812ac381dab246217754b560e5c14c8c7212b9e0deaa3f42d322af2a989784721a0db3e3a9105321fef9c4bace1669fd2c047c8aede016f8cd9aceceb5aabc;
endpackage
package dat_190;
integer pat_num = 190;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2be7e55cd16cfb23f2947fc4fe28f2ab33000218397202fd6861bf9f484a01626faa2ec0f2ce8fcc42a0f42bf6b22da560fbf8031de4178a1235c074af273d7b2f49c6b8db8b1745e500e52a36fbd5586542117b1c96920d3fa9aa69bb2dc7b9;
reg [511:0] golden_data = 512'h57003d9a565f0ca65d5dd9a90f1135e6fe7d0b082a5e0e2b4e0a2cbdb8705df241952a435946549cc088041f584ff4d27a536b36dfbfe48999339815a2f0b2a8;
endpackage
package dat_191;
integer pat_num = 191;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2b63694772e92205ad75c3cf9aace7d4d7bdde1030cc730710e4968faaef115a424e48e4ef48256b36b3c406add68061db2e5e18df2762339818f0a6c0dc209b493bb0d52d53b7f6ff6a480bcdde778ca63a40b86ca2e16dbc226ac8e0fe94a6;
reg [511:0] golden_data = 512'h41f459298d70197a922a4f8cb9f5f27dc3ede1dcf02d4052c411acd573a78fde74a4aea2ab7e33934194dcc38d20588937124c63fa666338d054299661a344bc;
endpackage
package dat_192;
integer pat_num = 192;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h62df28ab35ef638b7d545b4238162def8c5a8f9114f123dd743d2051feb32b1e4223932de39a96b7b06593d742ed47396f080614631ebaf976372fbb5bb74a0137eb1e2ce48ea8b6a09b0b066bf2d5afc9c76fe9ec32dbbb90280c1621df6738;
reg [511:0] golden_data = 512'h589945aedd5264a7e184069e80247e1932706562d0fddbf70a1552d0eec2524e103e4bee6841f9a10296f34af4ada77bec5959ed35307712b5e52a2458cea33e;
endpackage
package dat_193;
integer pat_num = 193;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7b0e41507469769023173c50df13eb6875d4cfdba697e5dab5bedff4720eb3e90fd9eb4a1002e1ae6c23f7613849b89491e50bfc1bb7c91a26eccbc26d2a48636934befb93cd1bee21e5f13bb272c9e4d10fb3734cf2b5e0c7a7db8fc49340fe;
reg [511:0] golden_data = 512'h689d8b0bbb4f902aa587e156932ef43d7ef0fffe820a64d749e988793b1bfc2436db74d7920d532ea7f6bc2e9018c827721d1b95471bba254d469930fdcc68a0;
endpackage
package dat_194;
integer pat_num = 194;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h560a0c20a7d3ac36df08729027a1bce4d89a5a47277f77b9b10d1271abf7a6d769c9740fcd8905fbbcf62d722ec935a3c6f1eefb6d7918cf7d5b0e7be211d9cc5812840a332117a9d3a31f01dc57c002ea549b85945c7cb303056f880e3d8c08;
reg [511:0] golden_data = 512'h75c2817688415d95fb5c5425ceee9420d5829ef2e567e273210bf3225cc06b0053ea50bac0b6566e81c8ed60e63cc9ba1f3ad9d415398c6c81b60c58a377ec4c;
endpackage
package dat_195;
integer pat_num = 195;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h217684c133165981d555e427a28e7b1f1a7b791a3e28027e6588f10eacd782814abbb27c46dd386cc7be3ba6f1cc7670dfbe8c2a8ff6a8b8fe6b0c20a0f98f00472cb9ba8b1aded3104eab5ccd3c41f552742ad528ff8c92d34483c604a5be9a;
reg [511:0] golden_data = 512'h1d7ff92b4bb58d95252639fd4c4044909bab589f3de88dc9533993585749e5ae4c7f670a2acb7ac03a0b8a706ac09705b614f4ea6966f9d4ebcb0771a5257200;
endpackage
package dat_196;
integer pat_num = 196;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h46fd4771d3979b06aa6f8c2aa69097e9a964da6e9e762094c7cf6961b1195b4436d4b377545b2d490731a0c198e7561347400e22d5c54f26928e759a1cae601168a1bb2c6c885d3b895f0230f3f3f735e41ab13c6143af4f5762e87351fd8505;
reg [511:0] golden_data = 512'h0e62c5cb2200380d3f319d43e9f3e654831b081937b9fc1f672b9be488d406687a1164cc76a74c619669533470c7a27f940d09b56ecd9c05d950a7ed74fc3bac;
endpackage
package dat_197;
integer pat_num = 197;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7f04b3c719bb3520d9d295600ac87d3e6007201df9711bce4530749e34a2c71a3f22b89c19b88ea2ad55494cfe29df7d9afeafc5c95c9c2d730c6d2c0083b4526aaa4238c7c18ce60dd101621df30af3f22b5e548893fa908280408a1b2b7f4f;
reg [511:0] golden_data = 512'h0a6b3985407e26195c821e97f7bd3d15e2bfe6438dd5cd1e27708e0bbeb76ce6330f79640ef6d47c94c51a48fba7d7c843064d4ba6e1336553ed2f88bb69522e;
endpackage
package dat_198;
integer pat_num = 198;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h73027ac511c9c807f17aadf03ccf6a247fd3d23eada9e8e61ec03ec22a8b2a9a21ad29d18a9326dfff5d4a066e810f975bcaabf709adf0dde319579d3b6bb175013d02debab3e30c97cf9f50844ba292f79084759401309d00379d6e2b6f46a6;
reg [511:0] golden_data = 512'h5a444bc21aed9edbb01b3ae9ba4aa2a1e114570f3cd05b8626bff12408bcd47c5c252354b41fccfa0b378c20374e46dbf68e23d9ec2598ad76fac03c5338f5b2;
endpackage
package dat_199;
integer pat_num = 199;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6251d87cca8e6e9824a3bad777dbeab7e4b9a52a0fc27f59a02a3dc8b8da6b15597d2c1caf74075df74a48356beebc3a415f195261356b4105df62909840895477fe6ea8bff20045aec7c5989b0cd8422ca5250f74f9555e01f4b9d0630c73e7;
reg [511:0] golden_data = 512'h43f3fc3397a3f36c0bb54043d865b1b83f12aa2436adb04e326a4e58bdf0b0da63d8c1b02ab94a6a2f2a8bd5050412b3e6209e54639d058b9d073288a60536fe;
endpackage
package dat_200;
integer pat_num = 200;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h405ca1be419c7699cac690c0f2b26a6d68933ed2e84056d875165767249ce0fb5a53f7bc77191a6ab80c486e649a2e70e78fd594487924e40e268ae061a33666264e57e22f6b06ee1f3f101d144a47b15478cc786950c896b768203fced72871;
reg [511:0] golden_data = 512'h75d92b88c3d9f691971c7ac3fa4d190233ac4927f537ade6d7e3f3ffd334b98a09925cae04e4d7b1e384ffb6f5f7c39f0121f9ce184bf6368b3d44c520d9734c;
endpackage
package dat_201;
integer pat_num = 201;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0559c5683d408fc4b086916561435d51b53a30ae036680f8c6f3397d270c2da85333debc3105641dbad5ff8f5377c793bad55df3d753d273642486dfa50eaade0a405cd50451dfb4f9a4334f76f247cb3a3e6dced91e95173e15979954240bef;
reg [511:0] golden_data = 512'h2bc263cba5427977fa6e17f813459a264a05d927a4827e85ac11e001efa7f80c1eca32adccd442d3d82bd62afbab89f916604b695688d4e638333cf35bb27868;
endpackage
package dat_202;
integer pat_num = 202;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h77c2d5f46f2fbcb235712e2192d70281170227c3f251529a21acedfe7496842373576dd64ebdea50587c30fc8984ab1c37eea0853ff2df99b24596509945793313ea34631c3164db71e71bb97a7d2e775a1cfa310ed92318ecf0c0a35e2189e0;
reg [511:0] golden_data = 512'h2a549e51a6bc4aa85a5e8f4f55f887a981891d0f4799990dafca290226c6a942551b3359bd7fe6fcef8973fa9211219372040cc261df8c8d1152f573c38da81c;
endpackage
package dat_203;
integer pat_num = 203;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0fc99be7cd0d19ad1ac3b5bc9b39f39e992f748df436c75eb789cf6dc257e154772822a835bd1645131835dc48010ec385ce139a79acbe7d0ec09a68760931ec027085ae94928cc12f56c55e23573a3c220304a6c6f6a333fdb8016336491d0c;
reg [511:0] golden_data = 512'h46329263844fdca3c7839fa9faebd00ad831f1580025d37716274ec93f31e09e04fa8dbbb9a1fe3c63ca751a2bdd6a14cb7e86e296893c2d21b1b361e97bec0a;
endpackage
package dat_204;
integer pat_num = 204;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4b0a34c5f9ce4c9c2e21f3b82215bd4e24b527c501cc363ca1a8ebda3521f1a13fe293bf449c0fee6cdc327b005271a6dd42d61768fe848ba56b9cb549d4ad4e713e9df7454650aa4125dcc7145a3b89154e499443be9d24d3a79e85adc73b54;
reg [511:0] golden_data = 512'h1259f1cbd34ff69a5647c84683033e2ba9f2e26eedbde09454165b0bbc5b46ee61d5a72a804db78a9067a414bfdf080204988dd5a306db791ab9636723f0765a;
endpackage
package dat_205;
integer pat_num = 205;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3331a6381bfed1c6dc4b774f01030825477bc22c72bde009fef7111cab84fdc5551774f20c7e69d9d4845ba00c59455fd28b69174ec54591c87e2a4779e2b098020319f8cc4f604cae2e74ba97bc8acc3e56a142fda975969e00445b66e17038;
reg [511:0] golden_data = 512'h48be6435724f0f69771d9a725bb27f850794f574e6e507e1f2e12888756c0ee668ba181a27e1470e524be314f7233d13cd58e71a1fc93a8358a2d9250ef9f30e;
endpackage
package dat_206;
integer pat_num = 206;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5be4cbf0193b9e3626697629959758db9f5727e3f91d779b81a78afd76e1fba55fbab8ac3bdd1f2d405cb38d9251ef4dcc08db537ad06c7e951a4ba1d82c67973cf118188cacad81896045c44a020ef6ef46931c5c05b31ccb47a0c364b742d5;
reg [511:0] golden_data = 512'h02651fdb494de24cd4b2c6ce814259bf4b9e353a8d4f6585072ff31d25da868408c3cb645525beb0a455a31fb0c75db998b274dffe66292062b6b372138398be;
endpackage
package dat_207;
integer pat_num = 207;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0a8f7ac76a3c44dcb7d89f0416851e57dde655ed4c313adce553f8b10b22ddb40b383748fd6d7954240baee3a78769f7a05771ee644ebc07825af4fc41ece1c85740cd38d556cef7c39016a3530c2ba51c1d402d72df22b835f19f92771f9cde;
reg [511:0] golden_data = 512'h680a21d21d694bc2ed96a1b83b914c622b10e3a9a0d7f290ea5fe2281ebefe3a77e5720be9769bfb1f01c0de30ae8e9f6983b585e25307dc9d53135b8b1cf97e;
endpackage
package dat_208;
integer pat_num = 208;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h21d4c251e1f74e8edec8bf2666de5b520c418eadaa1c0f2b94d000cc0b51c3f53beb79e1a6e048a2173abef3d8eeadcf8d4937a0b9c369685661a6624d1eab90336b403bfd98f8d652720d354b0c2701b3e0f48b7bfea01041943d3baa36ddf7;
reg [511:0] golden_data = 512'h3d1f4c37591e8bb3891e292be3bbacf3c89b29ad79f90f3c6602644f5ae8075a1301aa2296219de7910b65dffd402724656ccc18327b25f12ffa0308e23ba986;
endpackage
package dat_209;
integer pat_num = 209;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1344c3e7af4935cd409f20181c43e54e64fa3c04ae3a1d3f2ef6361392293d2c4c1024c8a88b6b0f4f19f66a04708ae8ed1c690dfc944e0c22dfcd41d243662b34a7ac95f9c15d190b132fe0543d37003aa156e0d450bda9ccaa9799b8b0c9b7;
reg [511:0] golden_data = 512'h1ad52fb076b93457c1cafaf58588a50fee1bb0efd1b81dd0f667df6f326c780e6ed9cab8f4e2bbbbd74a285a9d2155af172a40b00e6351a301c6b72aedfd21d2;
endpackage
package dat_210;
integer pat_num = 210;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h672cbc09068d0f6c8e9639fd7a9c6ac739a61aa5ebefa555baae4951c0677dea12e3cdb1232e43c6687a1c01564f46af46ad537a492e99f5a85ef6c5c183af62293b4cd8bb82c4098f217cb0623ce11fc931a8aa1bc8460562cec249c64e39b0;
reg [511:0] golden_data = 512'h194552c64f9ba583661646520934fa62bac9a5a8d4aec79e774b1f10ab0be2822292701e843fa65bd4d4843467c67206961feb45e2c46053855f48d81e7fb376;
endpackage
package dat_211;
integer pat_num = 211;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3d33eb8d4b5d58afea61d458a38693d2e003fc095373760600ed8eefa316f28b7af0715f7fb336c417c84f2f92481b01c04453a1771cfd8f996be9e66ca00ec95470e9781024dca1e6be480b782d64fe1213960985e648b2ec1c39216ffdbbaa;
reg [511:0] golden_data = 512'h1dc741cea512b6efec69d8d5ef40ffdb5b131d8fcb3228ecfc3a34c12e260bd80b3f4857ed18e5d34b7529492840f17abdfd52da975a6883b99b8b2984004de6;
endpackage
package dat_212;
integer pat_num = 212;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h18fd61d7a8cbd001b7426b90bf2a10a94ffcf0d36b0aeb28cb9f88922a4b7e7a7a0fdb59eaff17d68e1e3bfb85bc12e4b1ee31a507af836c32c325948c121f0a4a7dd192e2779605aa4456977f4c910eb39c4af98936c932f7639212c6e74285;
reg [511:0] golden_data = 512'h189532650078f2a2c23c3177006942961f90ec717fb2d7f69b4b917222bad5ee7f3f1b7735b6d8b95103f300f19d7f27cf0ef6496ae860be8bbcfc23237bbf10;
endpackage
package dat_213;
integer pat_num = 213;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4d31c94ed30b27ac10a7832d41b65fbce0f17e8fca0f0bf9686432bcf646dadf78af2bd4b4a91eb7773be5d5e649e8e9d642e43b7e3aa59bc4fadfdc97a7a5a009efe3a3e71a07e0a78338569b4bb627f28495b59cc58498b54b66c6ca64b55b;
reg [511:0] golden_data = 512'h4bfd7ee3a74320b0f3eb3b57f7d8dc778029c25a02ed3b9b9c8ddb40eea8c5e01bf45be4f8e0e951b4748896c43c5a4cc9f63b8283659e57737b62be6e3deb1a;
endpackage
package dat_214;
integer pat_num = 214;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h40a976ba0985f74097db165da61c335447157e4cb9bd09a9d46f132cb10265e64620698788e47ac6c2424dddc664a13209af56470596f93f10e28e6f28a2aa051fcd1996898766c53a9034dd131a80a1c2ca37e964371c203c38af8543bfe902;
reg [511:0] golden_data = 512'h5af8f4c60b702e579da619b8bdd6eea9e89874a6ffa52c64b7c4263d2c8244ba560d87dc1a72f6f95b718e28c33161b3ae3e0b53a96e358a7c9a9e89d905332c;
endpackage
package dat_215;
integer pat_num = 215;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0bd8b62eba708dec66e47b6954dca9d5a55d864ed051b76d6557814343c7401e40e8bd723ff4063cb1da7117c0abc9ba90f716df20f196020b49183b654c971278445c9ce58c51f91f9a14a2a0eee20a10612c43fa1d5c1302ad7e8b9f2364c7;
reg [511:0] golden_data = 512'h6c9c8b85646f6e5cb34eb0a5d56b8df3bd21677cd028193ccdc71bc7f31c82163ecae56cc4004084cfe318c9d5758887c07036c9a90d2cfbf8825a4fb83a910a;
endpackage
package dat_216;
integer pat_num = 216;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h14e1636718b1e48536dc85678e1538bcc19eb3cbe192fa4f398de6353af4ada24852e7593248134fb81a40bfcf724ec12f56c78b46b88bfaca0d47433bf9ee0a14bdaa68f761293074b5b09704cc6d5f383bd0af6b280814fe079db2910331f1;
reg [511:0] golden_data = 512'h78e7373689e0f5f4aa0e536356448dc56e32496834d89b5af04792f5828067722d9882ef96ee81511891f70974c8a5fdf778955b77a093fa7c229533d2723d94;
endpackage
package dat_217;
integer pat_num = 217;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h199aa42a458a7cd2f6e55f2cf49dff33a990c5ac5486998d214af2bf4472414e19c3657c508988514d04349cade63b403d91dc95ddd0a6b1b58a89319fcb4c4e3d2242a9ae8ab671461dbe985f935e301d27a205423e14cc347088ea86887913;
reg [511:0] golden_data = 512'h0e18f7477d8806705cbca879fdb6c512d7728b872c3edc7791008368d2eabca00f6a87449e978437bda1879a11bb97d3c8c65702ca732c0b75d3841ff9e8208c;
endpackage
package dat_218;
integer pat_num = 218;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h148ebdd8d805e773ec20a76a5ead533934889bc7c16861e785a82ae0c6796c3c66d062bae5c992c12d0bc88a761dc42ed47720441534f55bcb8fa76dc68e824e453a078dd8f51f87e6e966fdbe1caa4be509f626b81afb9d3390c0c36130f124;
reg [511:0] golden_data = 512'h7c3176f0a7707069be057bf6fddbc119d18c9cdcdf91b0a7a074b78e41da68ec4db222d57505941b7503a25bda24f5cce61325cc74a226d1e2e66c94ab2806f4;
endpackage
package dat_219;
integer pat_num = 219;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h45bc58bcb3f4aaf4c9c00da45ac89d6e6490e74ff6027427a92f45551602810a75bf1d8fd7fba7bb855b76e1dbe47656d4f4e4e1af52a77e294f91a24da3e8bf6aabca494309c4b77cbed5c083f55be2509d830058d506a41da9186e8464ecf9;
reg [511:0] golden_data = 512'h36d0c92868739fc43d41b3d7845db14f4c0237b796194ffff32373a3dc5daa2e777e57a01407695df87e51b78b6fbc7e3f8e9a697d4b15e30b4f07005cd312f4;
endpackage
package dat_220;
integer pat_num = 220;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h49264932456ed3e07770d830075047ac40e0fbd3e818de86da0e333ff6aa277e21d56e3dbe0407f6aa16cb9f09dce2787f8e9d7bf5dbee8ed54852cb25d073371fa9d3df5912014e9f95439b366d2ad1d380ff705c6040794b3a5317c912c20f;
reg [511:0] golden_data = 512'h39a2ba49eae79e4d853b0a3c9fb0d3d6df80d42730cdde3738dd60376511890c3cbaed6393107fa0bbeccbe9b8cb745d937a7a5e8b81a9d97db983a73735341e;
endpackage
package dat_221;
integer pat_num = 221;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h75bc24bdb42190deb5fbd4b8a1602652abdbbc311ea121ae1f24126a6a45cc2f16070fbbfa16627e6b358207c066239f81ad6e8ba3b98960717d75d1708b2a6f606e6cbf5b9e49fe351ac024f0896995f74c79a2859fb703b91ba428001bb690;
reg [511:0] golden_data = 512'h57e27c8fcd95e787a5649adff3eca783c8b2cf60ca216b8d112d336a4d13e9b663f1c2cc2b9863460c8f1624a77c5216391feaede49004220b469de21ef2fe36;
endpackage
package dat_222;
integer pat_num = 222;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0c17c196be116b956c3b4d6fe208a666896bc28ad50d8dbc2fe0f5911738c599580f5ccbc7e96bd43feafdc9ba7d1a4fb6f037adcad0325ffe2a749bd7b51aee0f77d07234aec777b4f824cad001bbff0694d79cda63010110b025a93029c351;
reg [511:0] golden_data = 512'h12e86658a92a2fe2c4b1c7cba99ca9f64ee7dc8801aaa125219bba9da49b1d62244ce34708f22a3bdc0e640d03d63723d088e3fbc8ac32da0ef3168d9bf403b6;
endpackage
package dat_223;
integer pat_num = 223;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h65fa73c7d6ff8d1c5da0b9c16aa12927b86d5bf603547bd677b82ad747d7ccbe30b28658fc1a9f2dc474ad1327215383e7d87cd0af77c06e4e2752e74c804e856a7e01836309d61aa2e596087a3634977a0ec825712664fb2dd7e6f25a61d9bb;
reg [511:0] golden_data = 512'h430e651b6526bf531f3aed00d0a761aed27a9038fa4fab4c7238441b65cdcbd80695974ae1502f265e80de09d865bdb4ff041ac4bf4c62f19c754197b7726904;
endpackage
package dat_224;
integer pat_num = 224;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7421e8d0921edc4d4e7246b85bb5edf7b0da0cd33f91cbddd3126798b75538d60ed0c0bc78069ad1e4ae4a09aa93f0f572c5496f0306631bba4ce56d5a8f5c997527ae360eec7e76157b63470ee42efd6aefbb8a2e903540e9a4361aaba8e0bc;
reg [511:0] golden_data = 512'h4247154e980c947680403f625603e72ffb246e5fd3a331b8f17335bd053a3c8c4ce2cf78d38ddf01b226bc3d274537cbd66f1f159a737e13a2fea9ca60389546;
endpackage
package dat_225;
integer pat_num = 225;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h147cade7f08842b2bfe5d51312a0f1db1692192408d14b25505a18c37e61631f1f6098209b525b0e4aa41749058f54a64205d56c8dd3963c55fd6ac2f577314f3ab9329ba242e8a4da4d8a3b16514c3e4c5794d60fde2a86859bfcde65c58c42;
reg [511:0] golden_data = 512'h1ebea82576eb0e77a75d61adb6ddac531ebee82e67b256dd3304669c5c4feb161a3e523fa11986fd5ae0959cb3fe06dcebd0c63cd095fc90f2c17cf778b7b386;
endpackage
package dat_226;
integer pat_num = 226;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5798523e35ffe15466e52741ba701bd5ba85e25aad201862bd07ac259a7d3d8322a8ba71e4b573a5fcf12f53b8ac9723b88899dfc4a789724d6def407dc40d7033c1645224ee93a3f6d8d3ebd59f6697b227ed9b5e5a46a60123760227fdebdd;
reg [511:0] golden_data = 512'h53bb66b3294630ee4e29b71ff3827c87cc3af5409b10e699cf1c55406bdb6bac0e0643a55035f3871dca5dc1db018617598bb825f9a5ee50c8a53d2ae632a9ee;
endpackage
package dat_227;
integer pat_num = 227;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h69b124213c0c78c8b8549309ee70fea430b404eecc1ce05e25a2332b47b60bd6192c03b10d6f3fe4bfe2b4615b955d01ab5084ce1372e6709d3f0a09d7f08cb922fc6e1818617dc4485a4342048a64c4721040307262b8124fec75eb15130ea4;
reg [511:0] golden_data = 512'h2ef969030c13659ee73ca3006ff036e6f8382a4612b6fc3341b0511170ffe5bc6ff2e074d1170f07ea75db51f1ec364d18d4ec386ea201707d51bff2d42054b8;
endpackage
package dat_228;
integer pat_num = 228;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h073f9cecdcd72d3acbb7c190ead83b22ea1535a5315052f278afbdce569f2cb612bfdb23b431f8ac8c473338602408d86aeb23a4eed7255e75872a48651d0fbc2c01a6277a80db6754be933a396399ff65b2f347f861c3760a0a8a2ce647e541;
reg [511:0] golden_data = 512'h09bce51a3b1c5383a0f76a385c2bd98b7a90ba84e7d0bca1db8a2371a0981808466f12834829b6a65cb5db840dd9b8c01d49bf903d1c3a40ace993c0215b25b8;
endpackage
package dat_229;
integer pat_num = 229;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h391dba45fa68e022138653aa690f214df75e36ef9cab25582ef97a0746306fc0664295f9ba96ff607133da9e2ce5ed5e36917ee8404804e6409ff309f84ef48922ad183ea9c7080d557892f96aec029106e738f0ecd37c0fce19f298381ac34b;
reg [511:0] golden_data = 512'h69b13dba3e7eedfa00836cffe9c3d16d5799a4a36f36668c287cc8695fbfcafe0ee4a68cc5a20acbf3381f2c039ebb7b74dc4b3aa9a2acaceb46908e46f571e8;
endpackage
package dat_230;
integer pat_num = 230;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4736ade3cbae534e40d936dda642a5634b3161e235eb45c8936c0e6f2436535520309298d18149b2774cd6cc404c237f7d25fca581220404ff55ba81e7af566019a53722fb42d9d598739b69721ef6d9e42b01111c69c9d427359cdb8b1eb1e1;
reg [511:0] golden_data = 512'h07f82adc75540171ca5bc877108c0dfbcd71d89e5bc0542a2694d581ef389b0473e0fbf089b3d18a67b364368752d3f440c3868ecb947641545c31d40586aca4;
endpackage
package dat_231;
integer pat_num = 231;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h06d2fcc0fd993cbcaa97d240276e86e08bef309487ee9c7cb395f69a0df4b1bb1654b459e4688fe38af1b9ab2ac122202f7590866388a2ab83b81f2010ddd43053279dddf08a0d8381d271e9370931e9699fbae01ffa8faa882fa17624d353fa;
reg [511:0] golden_data = 512'h4b55892321ca4ba004c7e88ceebe1e954cbad710e3dd2a686868211d7a01216c0ce10f1edc27c3a7b1525818f466ab74e5cca5eb7649852865caed5981a114c0;
endpackage
package dat_232;
integer pat_num = 232;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5721aeb721c6f6cfcdf1bae26b4c77e90a93efeb21cb40cac293b601e9e5cfe248926aa4e7301128c2873403d787ef2bc0ae34718af65cc5afcc105b621568fc6e6b069229c2c211c8c32c77e6b299fda9d026b5be5fc4f9b572eaf6b9bc5a71;
reg [511:0] golden_data = 512'h3cb0a047610f2f4c313a5945d0b5e7e03e4be81bc06d6a45c1c2fc8792f18c9a4fd366a8456fb132f490b7b071e6523230634adf75208e0accc14fd90624f6c4;
endpackage
package dat_233;
integer pat_num = 233;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6b422ca06e3cc5ed9169456cd5b1fb76f9dca59ca3784e01cfaaa9cc02afa04a7a74c7dfa9417a035ad4b588e71eb6ed00fea2b6721502c0b8379ac6df8b08a327555e06f31251e7afe56ef143027820ee38fbc5ffd772a94b06518f1effef09;
reg [511:0] golden_data = 512'h01f97181286d6d1c6806aa677ac3a687edf800eedcf1f95e6a9606d318d55c2233512cadd2a998a3dceadbee33afb4f75c97a4f86ea99fd0edb621120b8e712c;
endpackage
package dat_234;
integer pat_num = 234;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h67ff345d98b78c295604d6db37b1aeaf5fb798a04d7f3e839c6b42ccfccf425a31211b8cac53cefc3ffd2af677bacece15567272ff9e8c5d1cd9d72f52e3673e61e5b3aa1b3a3d9b2097c1c9aea003d16d1de7066e869077af3cafc75c6f55e3;
reg [511:0] golden_data = 512'h482d9efb61108c3cb3a7aabc5131c1502662e5a1cd429ba843bdfe7bb60ea6d26c7210c38706f5acf33fb35e2b67d9c190f230584c1877dd4563a8cc322248b8;
endpackage
package dat_235;
integer pat_num = 235;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h25dc0a8b589ccea2c1f6f90a5dadc9851a0b546793294c2a024d15e363fc77480180972ac167962007bb1dcff5c5ce0ec1b040a73659d77fa1b7668c80632b9d227b64b30fe7bde682bcafad3561a6a5f4e0e3235702fdfd01234cb310f9e4e2;
reg [511:0] golden_data = 512'h43fe29a768c095dce94a32c72de6ec310b1b3edc37c09065954f66be57d60726405aeec1dd38835ac3b3da0a231dd62eeed465d539f0282b79fcdd8f17961476;
endpackage
package dat_236;
integer pat_num = 236;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5e884987dc11a118a6c71341b81bfc7918934eaf74f0a9ebafcd13af1b4e015d37b41e3f251ec2c9ea5593b0b14ef7464d6eb0c78831edfd16443d50c31d082b0db6a82a06e66f9cd261f7905298d1df1ac13bb307cb567d6c24a7a43229a05b;
reg [511:0] golden_data = 512'h1c476b44611051db9636bf0f7d693343adc22196c342ae801bed274866119a242e14fb73b5d67daca662080dd05cca8b99b09f1dc7c240c15f502f96306803b4;
endpackage
package dat_237;
integer pat_num = 237;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4ee84fe739bba9cd7e80ff8b90ceef3c9c4570d88b1ef1090919f53d87f6326c34a3426bcc108b04f62fd215640ebf950eb708b74b3f1516c760aba00ed8b394779e08953c239727d2eebc61e4618705c73a3c97e2f1b4ee8d1ee5066b0b7012;
reg [511:0] golden_data = 512'h56f316a50669a2c4d536e0957efb866678c7a8d806279fd375d08b93a13d66e8423d42b0acb05b967450cfef65f639c411c05db274001cfbac095b7198144678;
endpackage
package dat_238;
integer pat_num = 238;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h43116608cf968dccd8b4dbf2894f0845073dbb223327a4cc57c0d7547cba50eb4542bd7581359be2cbe0acb2dc824d5a9540cd55b483cf68491fc82c94e9ce1003601946f65231e57331eff804c21121770068659595bcb57908fc564749753f;
reg [511:0] golden_data = 512'h6fa0775bd1974ae80670931ac5a81ac0bee41f6572a835c7f3469a6eb0739f2c2d090d543e5fb30af535849f8a51b0bfc27ef5b980b21ed42afa687c1c2a88b6;
endpackage
package dat_239;
integer pat_num = 239;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h05265ad01d73b2171433c687960f953ff73ad37ffab0f61e599454e50a52180c37bcd6f04f47db10a52884f199c6ac0707618db003627c1d8f2cae2cc589153c05b10e68bc5f39e87b5814ce2faa79ce398ec7d8cb077a9f8effa28761ff009b;
reg [511:0] golden_data = 512'h6663316eefe40e93101410ac2e7fb711d1f919007e4e7cf56632da49d34f66723784c467a82aef4478e125723129ee01f5f14212afffaf8826e8ee77ac535dfa;
endpackage
package dat_240;
integer pat_num = 240;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h63bff703959a9f9b7c744b97f3c1b579e735df9b29a58d5768c4ab2086189e7259525f51ba6e076e8d6da9c192e087785276cad832a6404cd43f30ffa2fd841a0fa5a7687c7d1eadff3a7db49b52d44e4fbe29248900c93f99493b759813d511;
reg [511:0] golden_data = 512'h2e4fcaf68c8609667d9bf26556bb8687b71d100939253a9f6b06d293b79fb0b8507838ebe0bbcb79ad35bf0cc3aa2dc3e1340708d7f3dc6aa6b40ee5502539d8;
endpackage
package dat_241;
integer pat_num = 241;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h542a295d5db345e776569dc640918683ff8e8a9dc43725dd832c244ccc6764cf39b42ca7b5ab2e798ee98fff9c9c5ec77ac6bba4d672f45374825f77ce67029e74e2e2c5c29fbc5d619caea0eb91b09c3bf9fd4c8107b6b9ef7025ae6190d9b4;
reg [511:0] golden_data = 512'h6ccdcba6fc40257bed6495da5b2fd75b55e58695db4f2cfdf30a0b06ccd191647bfe55e9a6946c7076985aa99d5bbe5cfc019487afe52374127fde96b6daa3f0;
endpackage
package dat_242;
integer pat_num = 242;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2b49070ef3cc23af3f03ef06c061def2896b083852e695935c0b5bbc654f454068fbdc09af6a520b558ac427aef1eb494e413648f0cb1fe828e01f18812f6a697fd21834308da6c53bcc9b84bbb1a842060bf868e8471675b015c5ac2a99aea2;
reg [511:0] golden_data = 512'h449e226ecfdde1ac1cc0d80545edc6e38da896b2a2032ac16ea2a9057137dfca6b6801b0522e07d7c568628333c4a51eca15e6ae4bf2d18fa767fc7ab223115c;
endpackage
package dat_243;
integer pat_num = 243;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h6fad03dbfdb7e5f871ef96c2fd7b177f25c21e7461420b192b865d93809f0df27dd639852a5ed81582c1c30067948298b001ec683529afda88e2c6cd5b8977bb2167dca454c694cb65d6eca9a0ffbfc93a5a018ce42948bf43a1e9d9e9cb6179;
reg [511:0] golden_data = 512'h6b663cbe8a076938704af4aead8eb3e2fc4705d8beb07a4a07a58596aeda9b62278676c465fc34af9f0482d7f92025ed43e0990dd205243ab1b0f7c4504cb094;
endpackage
package dat_244;
integer pat_num = 244;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7049a7e70e96d2a65780ed1dce5c4623a8fc596e8e7931e40435f37c52b53e8a75b9df9f4f32bd9acf2451c735b8c4c89ca6d1903119ce49ab8eef411943d2d3512bde4124ff8206ca6abc0c0581ba051dd4ef2acb2ec18824706d3bd9fefc34;
reg [511:0] golden_data = 512'h4f5dafbc02bb628eef5bf7ec4a3e9cf4d05ee8e363e92f82a7c9e8abcab4b9a23325ea167b09372442b6baa307f5ae5ae0e92c1bb7b8dc9c55ab5f3b5bd161ce;
endpackage
package dat_245;
integer pat_num = 245;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5894808daa1255466cdd8e38a5f63759b6a36bb946fa59528a2b6cc97113b46c49d0b2360e1a70c0ab9d551fa2ca8e3026adc242ee4aa5e9e4a827f365f8a64634a05d2e435b08989af0e76f86ecb051f172a74e796ed0f8f93f961ccd1fa63a;
reg [511:0] golden_data = 512'h15903e687bd5712b5361b692d7a9440a534f3f585c5fa59b1b6a6032f46a2b7c02067b0c131147a591af05d8d5c6400ff698ec9fafe09b41764a47a334986bca;
endpackage
package dat_246;
integer pat_num = 246;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7d4695794477f404aef5192c43709749edff0ead3ffd74a57bdf7be3884ea1603d5a6dae5bad2d5b053277f93214a89ac0efa7291be8885d4ade8670212d27fd3aabd30bdb38a8bc1fec964d4e6f6987ba4a0e5b7ef8df48099b39b47e04ced8;
reg [511:0] golden_data = 512'h329a164e382558d80295cdeae5c1d8368bd20eed3865156cb5878818fcb16940249bf8a8522c37c69f3fedf725f9327fd1fa0c66bc1ab676ccdaab53395ec6bc;
endpackage
package dat_247;
integer pat_num = 247;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4c9531c279b0812e2602e860293cda04d0a1487f81d93d37b28744a7c99056062caee051d7ec12b53863547e5ae44d337ab937c05a8b82693e942f3ffe5277a8656702c86bfc8d879868f5a521dd53a924cd8aea2dfbbb355dbe12e63417ec0e;
reg [511:0] golden_data = 512'h46bc6fd19ce74f9708e464800c018f1017bd5e5b18a399141795e662292be8004b30bec9fbef2f082327ce28876856c1cb89c60531b35228608a08c6a5e0c1d2;
endpackage
package dat_248;
integer pat_num = 248;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h592c549c3b863d8b733a14dd5926315daa3dc7bd26661039ce51354552bd8a8d0a6cc1c6162ecd4d51670e1d17dadd2ef57093343aa85e554a474d80a69e3e3e7e99433641db2ce85168181adb5aef04744747014a3a6d92ac447e28a441fc79;
reg [511:0] golden_data = 512'h0f0c2f6dadd440598cc1da63f8d38222bba145b4f6bfba6afb3d8ac5b110dae82bba2ecfec3b9072499dff3fa7b8f684d1d1cd03e61d3318dea68e7c2cc4e420;
endpackage
package dat_249;
integer pat_num = 249;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h02d980830fdbf9709fa15ce6a5ae70dde3cf1d57a470932c6b772d7aa629b9094e829a6e8d3263edf8df2cf819254a2efe449c08d07c6915f76d6549baa830e262faf636dbda96ca4c68aa794ec1c9298192dc679887550bdd95bd300201c5ff;
reg [511:0] golden_data = 512'h7cd91db604d8c35d77984ec669c43aa1e43caba5dbd2dfb77270ab5d48d27902155b0d830d2fffdfe3cfd022e7efe4a6b99f0018b5fae973942cc26daf0a7be6;
endpackage
package dat_250;
integer pat_num = 250;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h319cca63fce9b3db4a41615b6e1204d3cda99f29482c50d2b60497a72063c99f4aeae372b12a669beeb38593f4871a887316a5803f83714dbf25557f89eea5ec6086c343f0e944e61bda6e127d5a690e3ac4087c8d538dd2e2fef99cc3ca535e;
reg [511:0] golden_data = 512'h0cd2d45ea845272a40492601f2219d178e0446261517620336ad79ddc23bbfc2284eb696f4b12484a7f072d7dcdd6f5f67b2c5d56854d85e694f87cdc88d668a;
endpackage
package dat_251;
integer pat_num = 251;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h27a2e096eaacd23ba20e5b4982208733949e2b35a17f3b87def9d5626551d75e5ee80c3f62dc558840d4de3575f410f8eb22f8e12d26fd7e3d4021195004b2ae74ce020f4380caa3874e20e43cbb8a69801bc177304efd21d929754460e1f0ff;
reg [511:0] golden_data = 512'h0c7f136ef443772ae3f4d8c13e52ce71e290fcb8f44a6bbd21437d83cc36e7e857d464381dcd247832869e0a233393e96d228436b75068ba6c55f4f3bdb9bcb0;
endpackage
package dat_252;
integer pat_num = 252;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h434cd700dfd8ebc5219e53e55f5d2be9199ed06efed044f1d9ce0ec7e46e2c775157979494d0ebbd331fae77d33c720c878b17892540b13ac79a63426cb61c86038b10690a0d21804d09fecea68a6dc989b8eb2c0f9f42e6c0ca26588ecd08eb;
reg [511:0] golden_data = 512'h71992d49ea9a97bbdcff3c96fdeea598ad95171c32b14899519bca3d7f65350a500cf6d174d777d82c2b1f465b061a1632b92fc9e3bcc007b574cecb476a8656;
endpackage
package dat_253;
integer pat_num = 253;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0d6ee952552f7db979eac948a7a8ff98272e36c45b301df1ac1fcfac9db562fc62192ca9d8b38c25fe6daed022364d4a017219df2d62d9fa7e0e3a41be2750a137f5220f6461faed6d659d6beb73e98d9581808cc14405646943448c3f750800;
reg [511:0] golden_data = 512'h2bf3d06a58a65dbbdd32a2a627399d62d6ae1c147406ab9a1fecb44e3ad134fa5220b793e0a9bb1f0920fef6102019b2fe2e88295996dc0dd8195698d2f70b48;
endpackage
package dat_254;
integer pat_num = 254;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4ac1ca992d233e3b510a6f92f06750f4356475cb8199b0a9b2fba8cfb13721a8298829528d3f3739a43c6c3e56f35d81b182bb4cb741b12b007539de27a3078b7d2dca7e7c55fe8abcffb9734e6936c23129fb4aa838155427eacb14be7497df;
reg [511:0] golden_data = 512'h220b2f97ca80985f5bbf0bde2dfc04d78814dea62f7710b9357bec5a52419c7421fab873484362ab95d71362df3d625904bb8fce68902efda54a00daaa7f7318;
endpackage
package dat_255;
integer pat_num = 255;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3611b9f5e35fcd7e5460a0731df0605fe099cd85840af4d33dc0f0395bcea3d335dae78584bbeaf59e790aab70d333357d7092da50ceccb2d769f4e0d4bfdf971aa0c99b269706753fd2c0d210cf6a025bd721a5144902cde9a04e8d3d4820ab;
reg [511:0] golden_data = 512'h1c189eca065d3e3a5746a576ca55c3501b76e735268baa51e1be387741655c2e0e986e3d4302492a3be1ffb8c3fa0fb38ad9ed46198c133f309c547975326944;
endpackage
package dat_256;
integer pat_num = 256;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1e97000e6ef42c949f33821f7720ed6f63abf8be94057d65db4f43bcf41be13d3f4a23143a2a6f164c0f815e485b1c1a297ba51920acfbe556d993efbbd18d2e01c7ae6f33fb2ba6ac87f2627962c638ae78db2f2a7de8c7f091e5c5638054e6;
reg [511:0] golden_data = 512'h401bac5cfb72165585cb3ca1ebe2df072df085508a4f5aa33f48e51128add40e7c234b661f559ab82ae1966ae40f29b6d1df4e57b10d167e1aa1b5c9d62208f8;
endpackage
package dat_257;
integer pat_num = 257;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h61a91c761468f17a76d0f464e06f687d62657c4f711d3739a64d0813ecfb019e34fcb5134f846af1a5b334f07e09657f7f0d12f117f4ed1fbb9af4cc4e2cf679053e3a688372765d27713d7dcf2d11ad9ce8c222559baeda8d5ce26650bd430a;
reg [511:0] golden_data = 512'h2efaadf9b8c60801746f7cce85fc0412f5d1baef31187f4a0ec5779402c8e6ee4beb7695a8a31ec6b2c233f66e9acdf173909d0a79aabb4ac1ff4720276681e2;
endpackage
package dat_258;
integer pat_num = 258;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1f61c282f884f1f9059692c8db7466314e8aef6137f25aa3515450057e96a60e7326c4fcf98ef56f91aa2cc4c7b88a1cdc0ead4e4e502465052e93495a51f3ab4f918a4308c3cba431a6d6c6bd4ad1ee72001b6c1a5870f8fcb8f51d41159d79;
reg [511:0] golden_data = 512'h7155af39e90ee5ffa8a08f998ac7f95a75a7e6600d2a8adac1b1fd6beb565d6c3ad211eaa4a83187a83c9b8ccafea0fdb24ab796540827dfde78d2e9809d235e;
endpackage
package dat_259;
integer pat_num = 259;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2dd45306345a43c8bf38be5638f6d559b09f94c8ec97462b98fe4dd9c0e51a74450dbfeac61b5a8c86003a18730328f9487134036aeb03b2dd26426d19023b767a4c9efe31b3045733603f8d471c4834a8a21cd91c41aacbc584c32c710f18f3;
reg [511:0] golden_data = 512'h799639f3ccc92e5eee199921ddad422e856b7628853a8a9731bf0bbe6b639e8c73c72640a8e8cd42e6df742540981eb586b44d8a90a7fb78a62093f2d46ac824;
endpackage
package dat_260;
integer pat_num = 260;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5c7c3a8e0242fcef1ce1ebb535af0af6ee16ac9a347801eb9274bf4306ef2972534e0671cbca9951f21dbfc4a9c8885bc46462df5a9cd11d308c79d940fd75a13d88ad8ff6e0eca61f7087830f391a2523e0a00f88eb37f55725762473af2729;
reg [511:0] golden_data = 512'h1a724d248db1b6f3c0588bebd7318d52c240ba5a5518c58c1ae24d4aea4ef120086967a8c53cb6f196e165b66fe6a9dc9ce04cdca21406180c6bbdd8454fcfd4;
endpackage
package dat_261;
integer pat_num = 261;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0cf735278fe8cfee03a4e7979f5fb169b66606670ead026d8e9ab0ea47bcaaa56ef79100e9071425f4348ae5128caeb0af10eb8bd26631eec0b1ae38adbdaf5e0f0c32bceda829c93ffe5650cb2b4912bdac5129fc6195699f258f5bcd63b7c2;
reg [511:0] golden_data = 512'h319ebabddefb774d780e415248d6fd91cc72d76d91647e5b5fb4c6e6eeeff78c5d06ff505c418776806189035b25083a05a644fe18ba41414645fdbdc7456eea;
endpackage
package dat_262;
integer pat_num = 262;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h7e6dad4398fd2feb3cff0257bb404bc118193b96370caea050389a00049677802640c3af5d393c995c88410bcd414f03e3f8be0f3878e6dbc900f13fdb8229d01d6224afac8ed5ee5f800d5d96383385496a78f798ccfaad9b351ef59a4b0411;
reg [511:0] golden_data = 512'h5672d67972103072ca7e4b5314824233db3562d0dc25360ea1387732f58b546258cd07f461ced30a31542cb6112a6aa4aaa9de4ab397926d9e10de64ac1caab0;
endpackage
package dat_263;
integer pat_num = 263;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5b95b487d1c3ee1b379e0c38268a870d711ac3aac8318f82c66e99c9a35374d60089dcdf00f1fdb612bad3f0e122736856dda191a534ca6a6f76c9166e8cf3011024d34a7412784ae3588ade733ddefdcb5b39bc2632b8b324b48cea4f723e2f;
reg [511:0] golden_data = 512'h10b08f8d59eb1943df39152bd09f7a12392a242fad33ba8039b23dca1d63598033f29a83ad3793d488b1df7e86613537acb153a05afdbcdc71af1fea79e7256a;
endpackage
package dat_264;
integer pat_num = 264;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4efe13a86c66b82d5893ef1cc4b905453e226f89f145f5e3490ff7b872d225fe47aecd02446771f97190e6271908863e8c348f2b2b5a9c897fe1682f6fff0ad063c140c436c152294fd55cbbafa60529636befc675f4c76833d0d2e3537a5b36;
reg [511:0] golden_data = 512'h66c80319f25f2226235a0b084cee78e4c9ad9087daa5f73f6db1fc97571f3a263d7714eb0371f9d464d84c7017d621c6742032b46f3f98b479aea4fb72b0e9e8;
endpackage
package dat_265;
integer pat_num = 265;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h69e3683864f771df30f1e6a51ec56425bedaf045847602a15991767bb1b8f91f22e979f422cf5a7e1d75fc6e94a0b4f28c0de732e61429363b2c9e2d2aa5bef6123a65829d91ce1f8483799a4f803f94ae4e5f53193447b7b5c5f9732ee5cdcf;
reg [511:0] golden_data = 512'h180c3ecf64d35cae643610003d9e78a963b8ebca9204ad57c905bdca2dafad8867f3f1fce6b2183674a1da98e0570533b32b97c27887115e22754f0cc86143c8;
endpackage
package dat_266;
integer pat_num = 266;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5b916b035a9154bf653083a0cc7f5e8f528083e215706d55eae29063b99974263ce4c61138c91a4fe9d7752360410d2813902179e3e506d2e3ff02544e60dbba50204ba8c0dcd7d4f7813a1f8a76dd7eeb08728ab7f6ffadc31673bcaedef7ed;
reg [511:0] golden_data = 512'h623a4b613693e47100688ee250a44c5bdd3781e48acbc0be5d3c9e29a0dda8aa7ff65236cf08519dd5e8cb1736c2acad1bea0e9125093e56743cf34f4de40b02;
endpackage
package dat_267;
integer pat_num = 267;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h700f66b3338363ecbb2183cb4be6c19f9d23b912dc81c15f68d9b187cab5e13f3948cdff73b3d228d021d2c965dc1a7bb6b0a461f75196a3d9316721d2c7b9a75b65105686469b1ee0486549a050d90485652ce1e4a68438a75039f2e45b587b;
reg [511:0] golden_data = 512'h539678a3647885be3f17908d4900ac93675878efea79ce195a2fcdeddfdecaf07889f1592af73c73440b3f7f72116d0487657f835ab2264e2af3799ddc1b77ca;
endpackage
package dat_268;
integer pat_num = 268;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3a349204623bc4d2af881458cfd326429e08589447f32b72c0de7b99fb9ba7b560fcc33b73e359fe5e700f915c4453ed35d608d14b4c203edbe907edad996ba21fc7e746e627502a4daf14ab5d124899ea0404339b2227cd6f6f5a5e6a87e442;
reg [511:0] golden_data = 512'h22969d2c7e846c53487e7b828fc687d529ad4cb20a0fe41e9049a078118eeffa457db1b731c1052cf22d035602f36e2a93ebde3c717bdb05f4ebf1a0bef98b1a;
endpackage
package dat_269;
integer pat_num = 269;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h347212fcbb4b2a7c0b179d62ca3b9f771ec417ab29e2dc9792657a4162ea25ec1b7fb7c4afa69515b04fcb674e293f4c757cf9d1a7bdcc838fe871d2907e44a73b31e73b8bfa61834be786aab975a6fd38e9515a8fb4ca353d8db1aa94188a4f;
reg [511:0] golden_data = 512'h6a01f4a0ce27e703229e35ecf612e0cd03e0866acdd7c5b035b632124bf83a883994af661841c1a85304979c421ecc6a20701b4b7cfed504ac372fbf8bf7aa1a;
endpackage
package dat_270;
integer pat_num = 270;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1e0f18a4805c69ada32d8860616b1b2f62f56279463822ce28c5713ce89a2b737fa5484e12072cd1eea0260cb5f6d3119a18336a3d69c1824e8c32c60a0e3c663021869cdd5f88108483c89ae2164250e05b51e75e1167f8ccff670d009f3505;
reg [511:0] golden_data = 512'h05c78b068e925dcf2a5e10bb8841729a9a3d90f838aaaadeeba71c88694699d86a8d443f445308c881df7b13da47c8a74cb92a832797d511a1c1c13a3fb3a16a;
endpackage
package dat_271;
integer pat_num = 271;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h520b44f8b39084e4771943369f2a1edd45d4f9b813e6f13e6123dbbcb8ac81117150af8ce52ac8c4c496034ea88b625a6b658ea7fcb760aa9c1bde644465f2ba45da7184e5787e14aa824c78f0275ff9ca37973f32f9b0b5b20e8a9ac66f9012;
reg [511:0] golden_data = 512'h376651e58a52438c4653d298d97354e917c88133491fe335306dbc9a16d2bfc474e1013f9248f2368ada5befb3db12a69f9ff9f051cd85421d19e7f00a9e780a;
endpackage
package dat_272;
integer pat_num = 272;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h47c8a4287e97c0be257947d8c2cfaa13afde5d555cde7c11c1c1548ad3afd4b52ddddbe609bda22337b31ac76265973a38f0e7dc8650f1b41cc95d28caa5b19f38315001ffc9e14cf1397b5fd1d6644c8ff2e92c750db142c828d2c560f04010;
reg [511:0] golden_data = 512'h223e593cc0224b4e19f3d0e7ba1f67f777405623ac6e415f7df849ac0ab8a3e823bb79bd986c4c0335c40db2a734060ba95acb9dbfbff87858962b074cf07d38;
endpackage
package dat_273;
integer pat_num = 273;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0dcfe80762576244335e49991e1c047764aea37fee9def0859f9e993f2497ca3286b4361ff4a63a8f3ff44dcfa28fdd7102fe724be3187dcf52606d9f2269bc365d57a4a3a2fd8f568523fdd056ad21fc268368cd773b4fbb61ea28cc41863b6;
reg [511:0] golden_data = 512'h1961356ede66f7bd5c32fdaf6727896b1a6301fcbaca99140851950b59544a2609cc4da8e95d033303f5829b4fde247d685ae50a538e76c72d3dc4da9caf9220;
endpackage
package dat_274;
integer pat_num = 274;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h71def19261cc5dd3e88dedca97c8f91bb5eb91c43b5f1fcd78c7e0e3a0bc9c6b15f7de15b29437a856798d83e2b5e29f95603d5e7f541a40e6dd9b0c90f6fbf5702251206d157b0037ac655469640aac483d3d039b6c209849c88670f3d38789;
reg [511:0] golden_data = 512'h393f2098cf4bc40450f625c16260d13fbbe548209b768e5da0cb855803bf514655a8212dcb747119c26e4938a4a557841964acc3d98da36791debdd4affbda0a;
endpackage
package dat_275;
integer pat_num = 275;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3c630f2ed4007465e557607129f6922f54e67565d3bf373ea1087a96e3a7c5e67fa8cf56ee16f75e839f9298853605879f59b1eb9c5f28f3211f7fe9ed24dc37706225c98806cc489571edb00240f52888cf5c87f13b20da86fe709a9584615a;
reg [511:0] golden_data = 512'h1e4cb622c716895d27b3e1bf6efbdb380d449ab095a44a3b571416fe9ab6e6464d05777ba3d08f281adf9fa94407ed80cb8993d4fa4c3b1e244bd2f6dbbb9b76;
endpackage
package dat_276;
integer pat_num = 276;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h672f9668aa77847b4972e7278209b65945b5258959b2c17fbf33d7c1995b002726322c6b8d1a751833727ad647ee414405e079f96054f0190ee17221378c7cde332a6a726bd79ccdfd21e064a41d03536885563151e1a17275305c3a4de0a003;
reg [511:0] golden_data = 512'h18fb42739a6e348f4d394ce1b2f397c385bf60b878c7b3fc84b5ce98922ea952705c8a922d28e1500bb59df08967508422d05fa500da96f48d04a465461fd08e;
endpackage
package dat_277;
integer pat_num = 277;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h06aaa70e6638d809bed4c60be36ebbfd4f46cd4d2fbb01a85c47b75518292f3836d2f43a43fd14942dbe8d08a272857900024951271ac74b354e49c075d26a1a757a6b77c05570cc0c9508659da2683eceecedff8fdb8e9929351c6d43efde5e;
reg [511:0] golden_data = 512'h676f0baed9f19a085365cfcffa6c1e55af14370364fc75015b26ab27cb4b467a3a0e97ccc7b84eb9bd028a488c116ff20346f57cf89928057a8a443d935a004a;
endpackage
package dat_278;
integer pat_num = 278;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1fb188f2ab1b679a06822c16cab21325e2bb22faea08e6639b9ba1217e6a4e68708ac598c10efdfdc37e484de4c96d0006ee9bdbdf43567006489b0d6190e8ac2a3dac67d17606d7564d205f250e7ecfed2dd0978bab1d1f19daec91fc449a78;
reg [511:0] golden_data = 512'h6da63875dbbe85f751381f3f2b955bb0d0cacdf3e94d816b6282b5a7cb2425ea56a6ccd999ad0379fd3d0d64ed4eee808e61bff47d8f2348a17aa311a4999336;
endpackage
package dat_279;
integer pat_num = 279;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h2e5b3cd2ed08aff62be989f65c6b5ab063b80c423e4fbd0be3bcc25f2916156537dc85d6afa698bcc373e806c98ffe841dc7ad75abe5ad270e7360c9c14034a05bf98d90b76c40958c99d517b8aae26cec4d57ef421313a0c62d2bba44e997dc;
reg [511:0] golden_data = 512'h0df036dda0700ba833b8e28b7f4781cae1bcca37e0629137c5df10d0263ace0020333293499eea43c20df2b6dff0f772c5595980674750652fe8b3a14af92da0;
endpackage
package dat_280;
integer pat_num = 280;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h57df6ef3380a89a3658a46f320a9b06d517d8741eb09f86a67b88b70af86978f790434ae6367a9cfbf6c81ab954f14b9b98cc40c7b3c16394dac9041e64ed50e7b3dc55665765120c133c5d451c175899581faf38808beee5fba24ef1f797ba2;
reg [511:0] golden_data = 512'h511a5184452956c6891d2e66bd58ed8d30d304a2d380c9cb750952bb3277bbe81be3dbdf278d273df7bc0476bda543fdb827f43fd47d337ffd2f8bb03549c074;
endpackage
package dat_281;
integer pat_num = 281;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h55abaacfd3ed880ce93238aca18700c387e273f59d2351c3da2efcec119c2c5a3638efd5e1c15b6c3a98a5395164db44fe42c00d4fec0cd811be40febbafb459405b711ad806d8dfa13b1f89b569c720a43fad8242c15c9b95ee5d962c95f49a;
reg [511:0] golden_data = 512'h1b20a85420e04810d7e11f46b3fb9e17582c88fcb691f6a943c83c620031090036163dd947e4ae0358816f5ed66ff995ef28c851ced1e3126860e9c90340c48e;
endpackage
package dat_282;
integer pat_num = 282;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h76b9993bbf07f137ccd2d199de738adb83f84aa14f91985c6bbaa05084ab85a52140f71dc614b0a6a1d37fd599591c6a9c03c737bf0fdb9b9dc13c50465a67b35fbcc1d4a09bbb3431a97c4471dc98914a9d16b2dab142ffcf330b6b95756d14;
reg [511:0] golden_data = 512'h7b94356bbf7939d6de8e600a047f6671fa0834340ead054912419f1dd6e9313a36103aae14eb6fe2973a68134e651363ec2820b12df4bd052f2d1883bd421e3e;
endpackage
package dat_283;
integer pat_num = 283;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h476e203755c96b2066259f10e18f75934866d665e3031e88e5f964a07b41c44b396e27be203fa4d3f1861055059ad8d7cc353d51ca03e2eecec035bb38c7cd100a08e79cee9b1a5de04c8404fe4750f9fd678e29315f97d616a22b5952d2c1e6;
reg [511:0] golden_data = 512'h2567d9cf3afe5ac631cebb27111ddb4d7fc2a939cbf0ee94e8e985f4d9e5195c762fcde711d6aab9e0eee893cc5884f9a52027d332ef0c7af13652488ad2f6aa;
endpackage
package dat_284;
integer pat_num = 284;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h60ce9a2dae2570efbcd3cb34aad4bd49f7b477d1d0932046a52ca16cff2adffb39ebb239e164b1fb6a86df891b5d60433ea13ad75808d6464800591a9af87013039495270af73ef54b7063b0b6c015a91302d091296f0eb0fc48daf595a15df8;
reg [511:0] golden_data = 512'h6073f9ce67c0aa0e85a475ab871db34dfad09a791ed11f9851e08f07e5baa8984c7d5fc07be620233465587547657076daa12e44dadc970983f50609fb3e6a84;
endpackage
package dat_285;
integer pat_num = 285;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h4d879a9675fcca339b1ae78839953b9b5d0d343bcd382eec615b0901f47443e923e58569ee9f42404831c5998389a623c18c51c510fd90220451086d7ab415912fd0733e381a153bebf23ac5081d7706543eba4df863870c581340c0285a82b7;
reg [511:0] golden_data = 512'h432283b793117a11233ba90e49968c76a9d946ce320cbd10a4224eed7cf4078269062f76914033f865fbcd81bc3f0bbb085781220caf24b8d1d2782c2fa855f6;
endpackage
package dat_286;
integer pat_num = 286;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h250d32dcdaf9c137490bcd0b58cfee3959a8db9e916257dea2a5e6c59357c6d0532f93bf789526d48d404efa47424085182a99fa324164a166afb59f7a4fff1d0002f7f2114560dde01937d2af17c0be00656c9c3e51aa5bdefa15205e7eeac8;
reg [511:0] golden_data = 512'h73d0371bc2509acc9308a24a874c50ab1e224badeeec8edcd606c8eddef002e86f013f1336f8a7770f4ea847e517fba216b6e8f8a88109b7e37b25c4b75bf970;
endpackage
package dat_287;
integer pat_num = 287;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1e87278447507cd83d7022771745f246b5e7e36152047b5620bfe0083db8e5a07c179976adcb044d206fcd856966b21491fe5785af1e42567357a0f74acd017a7ad594e22244b53cf38ccb097f4060ba4ff923d4d3dac79ac353d182f1dbfccc;
reg [511:0] golden_data = 512'h523ce6ec0665368d11bc826a8f8b330717a85ca26ac153224450be0288b21a123a8bf5c4ba4c2737e0cd873bcb3fcba67203f9d9c27e9f89cbbfe4f0a7b37584;
endpackage
package dat_288;
integer pat_num = 288;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h70d13e43182242dbde6f5eab4882128c56220b62430661c39d1b8b47b2b86ea63569e39d5c92081fef511b14562545d1ae317293eceb7945d1dd810a4584013a059a5a016741add036511c0aa5f876165ef8cbb49f875f4e8451adc7a34366ef;
reg [511:0] golden_data = 512'h66e8408ad81ad5cd0f4d04a707e8650a0a7ca6919bcc0c6f4f2f4cd9e2e69dea6083fb84f8e662345a28ce96e749efec6cedd1a8820d596e44b39a202b041daa;
endpackage
package dat_289;
integer pat_num = 289;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h030676ac8336323be78bbe3ec22ce1a516f788e063b1fd357abee51dd006e56d6061ff62367b545f47c06eab5c3a3c78eaf94782c63c35e6b43452cbe1789f174cc1bdc431a2c5fbfa35ebb315bf857005e1b94a1493363795ca9b4f22769ca2;
reg [511:0] golden_data = 512'h582991c7d552741df2a416b8c65e3e400c3ac96d4ea4c8fe0c6058e8e934184a54bcdb56f9c9778a7ba286f76b674e62bb239d0b6d2ae20e142ebc33ab8035a2;
endpackage
package dat_290;
integer pat_num = 290;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3c6223257b877703e253cad686140a73f2239bf46e01d495227ca674ffb3438645c9e01d0053724e371c0545683eaa600b66bcec9dad550599fce43973b5e7e50c65a447ebece4dda1fbecaa5e7955eb5f4a0393167a23d6766f46fcbfcb1592;
reg [511:0] golden_data = 512'h1daf670e708a7bfc3159f50ba66c152920b0e927d851dadb599b60c51722547a575e596d32ded8b45d670a7193083ce2efba80e750ccd78c807e0f0d23c7feac;
endpackage
package dat_291;
integer pat_num = 291;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0fb90deffa2852e86e043911e65325448a062ebf31163d51558c65e66b4ecc4b269d31eaa569a23098eec49b67d6c7445ebfe3d39512855ddf899d0144066d08657a1d0174b56787df5bb53a202da741fb696e71091519ca0c5437f3d8be05a4;
reg [511:0] golden_data = 512'h69842be5abb347f14f1158feca5c356ab530e5cdb42b5828637068eb01ecb51e228c91e22c0eb2a488aec47a0e4c5e772ddf1f4aff339eb3f423f558c8d8d2d2;
endpackage
package dat_292;
integer pat_num = 292;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h17df916e8c3ff3f16d6a8b5e203ffc9d8db52824c4feb634295bb311f0cb16190efe69c27ebc976f369424dc909dc81eb1cdba99355bc2210e263e5aa76d8d1144f256c6d6c8ca0c439502237efd118d08ed0dc234b9f3bfff5b184564684b6e;
reg [511:0] golden_data = 512'h481e3b15a2f634d65bb6ae4c57f72f43ab4180dda3c3fcfb8881929b4f05d0e804996c6aa263570e9b9537f78550d722414999dcb833e92b6b42c607dbe6774e;
endpackage
package dat_293;
integer pat_num = 293;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h457bb8d7c5ccc7e90afd11f21296ce38ea869973e5ddf694254c013d29e24ea70475195c850ccbe22bf784a876f835f8d51ac4952be5a30b64587dc72809ee7e15c8ceaf7aff6cd63ecfe10b456f25416cee880321c53f7a6a5f38d7bbbd7eff;
reg [511:0] golden_data = 512'h567ac8fdcfb53b100e06dee3a4187b59fde1bc8205aa52d626fc4cc25d76906814164de052a4eddc1a1b6d0a6a1f12758d666c749e013c12a7e126ac84d8ad20;
endpackage
package dat_294;
integer pat_num = 294;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h3eee391bacafff16ec5571f5250c58a147f5e1fc9645e7e2b892d7b363ad43a5721edea6897e2897dfc0e37bea4a7613b8e29657ac0a750d9293a28f7457b700743f6af57ca7604db95c7cd6e94f4c379c495d5b6f0b58c23528e4ed8f96189b;
reg [511:0] golden_data = 512'h057db3140c6921a58c77c641400b5dd6ec9475872e4f427722beaf0bf81844c67fe64e58ea35efbc1b3d34e7da2cbbb7cae0daf75e55a6733c217b844e7e7eea;
endpackage
package dat_295;
integer pat_num = 295;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h10b8a67716ea68a94c81eb6a353f8b2e15e00dbc6895ddfc51085434030291bd67c239f90501e4a9c8e28d0839fa2fa887083a38232ab45c71be5416daf2b4ee70456adac48752eae03652cc8139b799ed84f951ab3ef44110bbc67883f2898c;
reg [511:0] golden_data = 512'h07f792c909217638ebf689c6f6035d222f736cdb40e0fe80b3f061bae464745e3d31fc6fb63b7a494f9af3db0d542d217478fa4dc7cb7c125818b3a614155a04;
endpackage
package dat_296;
integer pat_num = 296;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h0dffdb4f92c0772c33711f2980125484ee942f90416ac2fbf40ebd87d33671003d47959cb6d8541790b959e96e4bda2cbe5dd66b6ba049601708c582c3b02fab6c3cf585a8f5c8024ebc9c23a43bdf216b02e04bd2016d7ae5fbbe8e2664c2c5;
reg [511:0] golden_data = 512'h5e4216462ec38a09b09de2639992145fa49415bb5a3f15a11b9254ae5b18d5ea5c7b91adfe30c7db1672ddace567e2b03a13360978a8dfa328300cfbc23afe66;
endpackage
package dat_297;
integer pat_num = 297;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h708ac65f2c538521c1cf43b53eadf1f5df27a63673a0dafb3e345c203908eb9b31837b0255ba317ebdc5730740d94bbcefd5537138b85301f7a84495bf79f2050254de82ea3a71838b164742d9dbda9b6a9910fa008109453ea043f146ad7d76;
reg [511:0] golden_data = 512'h78c4ab62f4e6028a7172b83f6899a73dbe205327350da2dbd547d145adce8cbc0a3e60198af50811eb627c34c777023b8c991e64311a004fcc322be2c6631664;
endpackage
package dat_298;
integer pat_num = 298;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h1c7a71e8fe76ce19d7933188fdb2d91d34e61b1aa556812f16b8ecb37bfdb5cf297850d219afd53ffeeb6ce77c91ec10e1896eca47c969190b0bd5a50236f97143eeb031003be0aad49089c6f9c0a67101abf007eb1c7036c944f1f7c297760b;
reg [511:0] golden_data = 512'h449513d4242b1dd472626770548a425e0997c2a8ed8c9e901b8984d483eb82ec4f4f97c097a59095e2550351cf4f21711dfbbaedbdf794b5009c4b2e8098e688;
endpackage
package dat_299;
integer pat_num = 299;
// M: extract scalar, X: extract X-coord, Y: extract Y-coord
reg [767:0] input_data  = 768'h5881eee47b618ee3c5fc90c4e31e88974b5c4d246fc5dcc658ae41321e514352698920076b905644ec8177fb5cd2ffa510d93ee100982d3f62ef07c74927a17d447d4d28275dc481d2ec3af56c5c4c02bb149a3fdff689f8848ad3c69d3cabbf;
reg [511:0] golden_data = 512'h5346a81cec990aa7ca1939764f06614f3149dd0c376aaddd8678aec49325611e461eeac7aa634705e162a13e737a6aa56831d59b584e35e07a9976ff47d6e824;
endpackage
