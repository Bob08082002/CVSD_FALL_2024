package dat_0;
integer pat_num = 0;
reg [767:0] input_data  = 768'h259f4329e6f4590b9a164106cf6a659eb4862b21fb97d43588561712e8e5216a0fa4d2a95dafe3275eaf3ba907dbb1da819aba3927450d7399a270ce660d2fae2f0fe2678dedf6671e055f1a557233b324f44fb8be4afe607e5541eb11b0bea2;
reg [511:0] golden_data = 512'h47f6a5d15e1a09495f9216eba5253538db62c06ad333adbcc86932c069f00d26465032bc1d1cace745d1b3bad5ca1115805ab1512361151d1c84c68aa2f54468;
endpackage

package dat_1;
integer pat_num = 1;
reg [767:0] input_data  = 768'h17e0aa3c03983ca8ea7e9d498c778ea6eb2083e6ce164dba0ff18e0242af9fc32e2c9fbf00b87ab7cde15119d1c5b09aa9743b5c6fb96ec59dbf2f30209b133c116943db82ba4a31f240994b14a091fb55cc6edd19658a06d5f4c5805730c232;
reg [511:0] golden_data = 512'h7a3afed80c2ab24733d7a3cf8b33efcd547e88fabc71b39da58b42a26e6c606c6cbfdc595891983cc17335e1ecfbd786b92805efbd5be956a142f23285f29f8c;
endpackage

package dat_2;
integer pat_num = 2;
reg [767:0] input_data  = 768'h1759edc372ae22448b0163c1cd9d2b7d247a8333f7b0b7d2cda8056c3d15eef75b90ea17eaf962ef96588677a54b09c016ad982c842efa107c078796f88449a86a210d43f514ec3c7a8e677567ad835b5c2e4bc5dd3480e135708e41b42c0ac6;
reg [511:0] golden_data = 512'h668e7ea762ae11fb5159d50df7f92ee488c0f5ac4266701687de38e61cc5c8062bc1a2c8137938914f9b6e42763026845c6ee2c134819c7ba755a513d05c6ec8;
endpackage

package dat_3;
integer pat_num = 3;
reg [767:0] input_data  = 768'h58c56e7173256312a6fa3a64c48d5c487f9fd281cfd4dc3a8d8479fa7f504e086dee2e8e0a13f5034e2b3f22b8360893b1f7e7565c6e2e22a64131960f6cc2c0353d4e59a1403502e9644c3d40a9af324c3f24970468cc8433e9617f09a1f13e;
reg [511:0] golden_data = 512'h2fb00f496f8f1ed97383758f53375643a2aebfe60ace4edcb165b0ccd7e3e8e410d9f25795e9873de3ffea0edfac077b7a09d1afa4c097d57f62672a781a9ef8;
endpackage

package dat_4;
integer pat_num = 4;
reg [767:0] input_data  = 768'h75a00db83aa922f506fd567677800dc2a691eb091e650327233f5cf51ffd2f9f1afdd93edab4a216fcbe9f5b565a2154e725fe65400e653cd2ed9cfa8857467025badd6d3bfb7912c4d967cd2cb67c11fa684d8cee461812ad832410ad50972e;
reg [511:0] golden_data = 512'h299c8b081c1bb7661d23332826297140ead0348203f863d187052a9fdb9a3a521c15873a90ada577f4ea8ee86fd3d9c7dcbe8318b3a87b81847548ad160183e6;
endpackage

package dat_5;
integer pat_num = 5;
reg [767:0] input_data  = 768'h6920440a5b239a3d46c54d4fb26de9d4d4971c34c11248cd2e5a984ab5fc957d49d45f119c24551b4c10659bb0ff7fcd4e6ff685e4a253ab0c7104177276dfa242cf1dda8512a43c92fbef5dd23da28ba99faf3e9248751b13a7c763f11fadae;
reg [511:0] golden_data = 512'h1c7f61bd0586f794aef978927f93965ab01f1a4239663cfd2d6361a5b41463b05ad679c25fc48c36e92caffcc66314a3088faee43e53521de31568aa398383f2;
endpackage

package dat_6;
integer pat_num = 6;
reg [767:0] input_data  = 768'h55023b21c8f640ee5dcbc9204e9d1d12e8e740dd612cb38e6831a86efa63df996e7aa3b5ea917c904016e8c6c9639abfabd1371262548974b852064da51db1fc0cf4fac308fb419900617c9d54bc87511af300b8d165981e8cff7028a63ce1ae;
reg [511:0] golden_data = 512'h3ab421fea71ca2462faf1f225b6e2eb90a8f84d5d3c87848f8b483950ceb6b485a4eb4d890852b80ead87b7a19c9d2bc6f20e2ce907244a9af44c9654a1aefc2;
endpackage

package dat_7;
integer pat_num = 7;
reg [767:0] input_data  = 768'h4520c1a98bfd08b6fd5a73ae9ad57fce8c159793772b288e308e541d2eeec75f23d41ae8f087b179aef696bd675caaff32c1f9fedb62063a81ea2e06a2dfab284b0846a32fc2f839dfb3dfe3b453174aa76e66779da463002c927ae07f2701b0;
reg [511:0] golden_data = 512'h1e0100e2e6c6f972af2f8b1de3229002850bb693dbd873ceff042ef7009e27602821e0c60abb5edfd2516d75572c929973b5939849b10d6c6497770bd1959c64;
endpackage

package dat_8;
integer pat_num = 8;
reg [767:0] input_data  = 768'h3edaadfd218f9c25b4b26f2fad9d798994888ae12084292f08db1a018c725f881aea85224d3688f536cfa04a6ef7d58068aaaeceadb5f016046c5832fbfb7e2201bbde401eb60c52bb5e82604cad725b2f5ad3fd8f9622954938bbaf4b0396ac;
reg [511:0] golden_data = 512'h3fee452b0c385fbf0f42b373e3e0f51a12f5bc94b0b128f9c791a0d6164654403924554bb9985994139d999d65af9db5358abe088223be5f92b965751a5a1282;
endpackage

package dat_9;
integer pat_num = 9;
reg [767:0] input_data  = 768'h5521019add4ca443961d0e4f3c0f3c426f82cbf69c31e36bd48546162ff2e78f31162205421ba5a68dec939e24fbb6c6fd99c70aa040b3ff347eeb8525461dba18370b68eda97e4e672c82b0fa5c40acd2bd672a4e140b110bef812b383c9ae4;
reg [511:0] golden_data = 512'h6b93b232e3d2b36f266f31af7d39c1053dc5942edf5ea8ca0df65f999d94469c57154f4a640ab0943d64d00ce8500ca779942d6da479fb4dd53bb3e67f9a99a8;
endpackage

package dat_10;
integer pat_num = 10;
reg [767:0] input_data  = 768'h24fffa968105ece7d927a5a90b0ffa8eaa69fae0cb20814828e720e96d175c9d7ebc7f1be8ee62fb50678a9f4c9608e9f6633b2890ca0f307c488bfef02fa3783ef5efa19e1cd18aff98ef21e6da3294a48f66699a51cc66d5c57b4595d09478;
reg [511:0] golden_data = 512'h5243d3909e38a265492bb4ec37872a67f4d541c4009dc9ccd8ecebdb1ecfb78c5f68f3d07b0240b79eb79b2604c518b0181303f1a3a7c1d7a7450183e56f4c5c;
endpackage

package dat_11;
integer pat_num = 11;
reg [767:0] input_data  = 768'h590ee8dd33541cb4f0fb9e546a6793a043155acaf5c6e6425ba4be3fe8ffb4a243f949039a03c559c870b6e0a892c29b0c3b7d0204462e8c53c116598374aea0780510bbb026c0a35d6593fb903f39e7c791880978f23932f4e3490814eed7b4;
reg [511:0] golden_data = 512'h4d1e84521064c4df57b3de547e6be78fa7161f5583f3d2c2df58d051b26042127c9c909c84c6230a3c3d2945468d8afbae31d2606074b0c22e550b6ffd0d87da;
endpackage

package dat_12;
integer pat_num = 12;
reg [767:0] input_data  = 768'h45ee9758068823547aa0dee25ab018af52187ad09fa5084d050b28690a03684153349fcc4b78374780d19222bcb333a51544a6667d04fb95c0b4cc7d4efd96a0616a8aec4ba8f060ca7c9299ab455562502d1318978265a72dbb0d6542610ab8;
reg [511:0] golden_data = 512'h3a36d43aaf44e378deabc790108bcf49dab98c693b1ec51053917d445fb0db962785113dbd01a68d1ffcee1592993b2642d5b676fd5f564cd99a0dd915cfe332;
endpackage

package dat_13;
integer pat_num = 13;
reg [767:0] input_data  = 768'h20ebcb58c602d7e6d7fd20422307d3d1bc388aa7404b055a0a8f81b50f0baeab7b23c7e5da7ce6f41681db224caa6269ce5cf30f2c5ba116c79b62831acd22866e8267b9762568ef7a4f74ec44858bcd8397bc3fd5d6c07e8553b1442b9c9ffc;
reg [511:0] golden_data = 512'h442a537100af1c26b4e424e3c53c421083c7c8d3ec179c6bf0b498bcb9e38e502adaa6e00a35262ec40dd9c19a40dd6c5a4b88ee684ec37cb1fe1f9a5ae28eae;
endpackage

package dat_14;
integer pat_num = 14;
reg [767:0] input_data  = 768'h1d42b00466a7799de392edec7f712adf0b75e8a81910f498e0d8cf0e98d3af41039370abeb0f739d35a0788abb944eef7455cdaa77889ae2eeb334a2baeb9ff81902bc6553576f2e55dfcc833d2501ccf89b18e640a73bee84a3af5a3c7d41c8;
reg [511:0] golden_data = 512'h66e51481459649ce3f3ae57ad924f0dd22e4beba2c4028b19a26a85b45bea0686999ba4a3a62af50c19f5345ffcd8a2d169d3369f079a410e55ab6770a09786c;
endpackage

package dat_15;
integer pat_num = 15;
reg [767:0] input_data  = 768'h1c8bc355076165f0d3e1d7b8ebe213a4733342e92c03406d8f05d8efdfb35ce81e182637db3e36e66ba14ea434d99f1bb6eec588de2c489661fdf96b79065d040124f976124401cd891ef3ba76074bee8171583f3a60c6988dd71ca77632469a;
reg [511:0] golden_data = 512'h1bd075a86b87fd2fa51d5d5f46339c1a190df05fc05b89d41d3c749651d000b076a3593649b75ff78c705c56352f0b4ac4a4dcf932712c9339c4e486a324a8dc;
endpackage

package dat_16;
integer pat_num = 16;
reg [767:0] input_data  = 768'h3208b749f0d73df295465417bf0ef085672afa9fb1fd0e720d92c3a42e4af7286a12da16cbb52f989c24a1152f68f01fdbb6412db8546e096ae38adec2be4cb21b2d77cd95b972e6a48dddb7f37fcbf67dff7b8370bd3c980e940ae9e4da3f90;
reg [511:0] golden_data = 512'h5e00f491eb44a48fbeea1a20dc99f778a9bb1d446414d18886983fb76d8636565350b95a94557443e0816bd37cf1ba7e27cc1eef5197bd37f3f3b94e80222914;
endpackage

package dat_17;
integer pat_num = 17;
reg [767:0] input_data  = 768'h11b79663a6dc632d8d4f359e16180a166369550c9a54ef659df3afcef6ccc32a60acd118ba7beedea4afd3c5468e23012761e074363103475fdaf3958324ce544724012f419a6aa37d24f8abc2f0b1cb9b2350b37e81b9574d16d84450cc7374;
reg [511:0] golden_data = 512'h6e9b18f5a0ed4e3d67d9683310f6e03583009490d01a84e029a152e44b50b1206e3c706494406daa395c01f475c0b6cce57b6eb1941d11a64aaf41c9dd8f3458;
endpackage

package dat_18;
integer pat_num = 18;
reg [767:0] input_data  = 768'h0f04b0cff169779d8e0f65efe31af4db188599448623ebf962238977d5096e2f48cf5b0cc2665c46c01a84f593692fddf5aa578326d639bfd90296a233d505920ae45d47de6e516992faa309a443ffdcd51680c45d46c9a03e65b253c4654a5a;
reg [511:0] golden_data = 512'h5bbdd32753b3ed4238f3db5074287f14d4b31a43b862d41980bad8d0cbfc69cc32cdb49ed5f568391443d5c64c2ca395608fcdaef7a0d7c8f754558e5afa7680;
endpackage

package dat_19;
integer pat_num = 19;
reg [767:0] input_data  = 768'h082fa84e7a513047d3caa86116dcb08ea4a7d22b3ca17ce6da33f3b856288c703114b9dcfa667dce9cccd38d89123c65528994d0bcd368a19c0ca60009eb0c44401b3ec8d4205390a56493b45c29bb7babebfedf3bca74e1d920edb523bbdaf0;
reg [511:0] golden_data = 512'h5d589f3264d09a56534dd9707f13df0713400d906d78e3aa4223009323301d38157f9a091e5e1e3f5f7968560bb1d85e4be53a72263691e41cd8a7ea69151d0e;
endpackage

package dat_20;
integer pat_num = 20;
reg [767:0] input_data  = 768'h355cafb07df68025d6c6d96e84b56d3543399f5dfbb97c2867c1e4b640f8c1f6120b0d4efa6ae60666571dd765640ae5ee7919ba7f0e2963579d3b1296f5e07429deef8b903334654b51a8d40a20a4024afe13534a6cea1a4642bf59bc7790ae;
reg [511:0] golden_data = 512'h2601417b9c9bb5cb739a11b4266ab560d29fa603a2b5445ea7bafad47e0eb0a6471c8abb23651caf796ad521554d187b4dff1a99aff300cdc8b7012a50bb3498;
endpackage

package dat_21;
integer pat_num = 21;
reg [767:0] input_data  = 768'h048e33afecc26003f21cedce4f8bbc1c58563037073e17cfe6d851c124ba431b67339aa4f744b2ddccffcd2b49027babe8716eb524c4a8b5b144441935cd8ba635a15e2ac8af9d44cbab63a932ccd845383b13147c661f9551bba0006662c9e4;
reg [511:0] golden_data = 512'h0b50041eecd16f165947336a5a8d1c57e67119e481f3ea8d307aed9c1661c0b61be5825784c871d519dfe842195c046eebb22b7db45886dd2b9263597790b934;
endpackage

package dat_22;
integer pat_num = 22;
reg [767:0] input_data  = 768'h0f7e9c7f2075dd4794bc1844487d4e1bae911445e1b7aae21a6bee5bcfd56402457b8114733a4abb91985fa63b9f04cb48ec56c1476ea0ccfbffd90e0f2c9d2c1d1993ccac306527d270d31ba0e0a7465bb8682725dd3dcf28e5b9e42c0f3580;
reg [511:0] golden_data = 512'h6deebec6c68d57429a3bc1e686585892f554bed3084ea9feebfc771ee5b2642a0b68d37bc17072b1660bd46fb9d77d5cf48d9b2348d8de7fcad74bf218902312;
endpackage

package dat_23;
integer pat_num = 23;
reg [767:0] input_data  = 768'h7eb8993d6c91a2a9ef11a26d1635ff72136f77432b3dec24e2af18725872c7f37dba9915d57d7c38a7f43c6a5f1d54fcd3e2ef9d16936f29068c54418682ac3e25c40e9c52c8df5405244da6f133aae8526aecf4279c7500eef0022949c225ba;
reg [511:0] golden_data = 512'h31c181ac8bb3e7d1468fb05edb34f75d204e96c85c959c75aa415dffa8066c906e304b5b0bcf934a93696772d6c7fcd988ef440467dd14dfe8fd092f7d43430e;
endpackage

package dat_24;
integer pat_num = 24;
reg [767:0] input_data  = 768'h0a3db750de6fe0550df297d4b8cdd092b054a50a018d8ebb758ee7aae73693f5102ef7e276ef9ab834458b71a8ea12443f1477cd776a0efaebbfa0f5d1f7af3c5c48b9bb22f435e7944fcd9143ec7b63ca62c872ab0a9fb3c3eab76e1c21b258;
reg [511:0] golden_data = 512'h16117483aec7d770f657a0bd6c1ad83692653aefccf5cb6e735d774c57bec8ae75a5a2dee485c9611e495d87392102f8d3c83dd9b01a7ed1e1552769aa10fa9e;
endpackage

package dat_25;
integer pat_num = 25;
reg [767:0] input_data  = 768'h61ace1265ce96258c9564e94b45a2d45fdea38c28377725776135112ad7972ed6a5a2bc411d04917cc35bfde1174fe62d70232233231853815ad2078367bf0a01dd491542d440b00fc5b8c87804701a6f6daf9d79d614432e3bc766be65a7c42;
reg [511:0] golden_data = 512'h3d816175bc7d4c75bd86960bfc2a7a5e8a40b7a98bcb4c0f0eef8d6c3255cbf83ed4f6cce7b6b0956f87e0dbf2edc3506b141020f116d6812d9212ccaf3b7de8;
endpackage

package dat_26;
integer pat_num = 26;
reg [767:0] input_data  = 768'h575454b7887b02a72ac1759b8910cdc7b19ff1b2b2aff5df23d065147324a661453396c596aa18499104da10c7bc80de7d355b1513dcad6b7703ab413c6d042e6150f9324b461f7cb42006e19bbf2ecc22f259af0057f1dac9abaeaadc9cc130;
reg [511:0] golden_data = 512'h1abf95e38176aee70ab8e07bd56ec514ee51058bc6bb6b81ce095697e7decea442e329f206337faea01517ec8fd3c42bb0590dcac29e9f53decdb05661c317a6;
endpackage

package dat_27;
integer pat_num = 27;
reg [767:0] input_data  = 768'h0daaedfde5061333eae65d89119f779b5528699a31cd4137436a64bad2976cfd213db9ecaebc667949ab6e5931d09c53d403e7b2476b76c72099911d50d9c986438f04b57cb52f4490c09715ee86a8373aaaa014731877d8d998c7c198f08fb6;
reg [511:0] golden_data = 512'h5de4ecc4a5209115ad6ba6862219db7783a4b18e20e1c1301d9337049c11ff2022de266a05e43e31700bdfb8e2f56d3fac5509ce02ab4640de3d58391871dcf2;
endpackage

package dat_28;
integer pat_num = 28;
reg [767:0] input_data  = 768'h05544f77bf01753104d92679f020a777a13214d430ed2bfc52a841c8d1e6f2e35352ad845a1d5c3624c495a053f0147be9bfb7b2531a8e5965806663e8bebbc40883955e00b8313eed47ead193b6eed4dcc6f73c6ba10c44b14989db2806caa2;
reg [511:0] golden_data = 512'h555c5350e16e0a93ab7b8726f51fec487855ab2b8a23d21558a6ab9f0f4629d25c2361d752b7f3708f2a13eee6da3f9bf00d92deb48f8d9bf488573e516e7146;
endpackage

package dat_29;
integer pat_num = 29;
reg [767:0] input_data  = 768'h56450a47b343021bb4eb2854acba90c176e31f94633dc4a4786e48967a8c31925efc2edfe826762dcbb37c95f02524dd3aab6cb85b39c08b1c5de67c0ed6940a6b34303374306fed24c2d0e2aac3ee83dadb2a19c49a876c6cb954b8608692fa;
reg [511:0] golden_data = 512'h1fa65f495011b23e26a272b9630ea9492a1f26d2f9e36a2331d8d3e1a465c4042c27bd31f4a23b5ad111333bc098d8843d05a3d52ad6284f9cfa6356b6b4959a;
endpackage

package dat_30;
integer pat_num = 30;
reg [767:0] input_data  = 768'h787d960ecccda4f6343bd91d8cbdfbdd89af63a59720b64026d8b2f430d49da400bdb7d786d3ab844ed3334845124ba142d8b3f9d8d3dd80b85f7194bd5fc5827ba9c49f066caa86d64172fb8104aa590ccdd55edd2f3c4b75fb64e31af64bc6;
reg [511:0] golden_data = 512'h48043806f8858a015e7b09adc68441de6a67fa51701052f8ebca07f1f3fbe7220568469eedc0ac24209ebfa23efedae28fe840f570251185be6d1b9977ba9262;
endpackage

package dat_31;
integer pat_num = 31;
reg [767:0] input_data  = 768'h312806a6aa2f07e642f0fe5d207c3d659b8bebc0aed511f0b9a4da88a806e3ec6c0f531b56d936df0e908610b8faa1c65298409ba6f1a7c4bce2a98e6152d7f22a998e431855d18d882724d58c4c7dda4efa7d8880584244b0087beef4f7180c;
reg [511:0] golden_data = 512'h29f4ddbaccaf4f69c70d79ce848c7921c502361e3aa0eb0397c553c2828b0b1615cc80aa8c72a3dbfb4c91388c22c199cc3a8f8b9fc98e896aaae2e87230eeb6;
endpackage

package dat_32;
integer pat_num = 32;
reg [767:0] input_data  = 768'h2c7b250b870192606e5532bf2b0e1dcb4073bcea8698b560f60f465be2ce45602f6745a3fb4659d020fa932615a9baf279094085c1fde667e3005e3bcb88f0bc1bf4c5d2ce19fc999c9396d4c888ea868c89409344dc1296ab933e3aaa9e33c0;
reg [511:0] golden_data = 512'h3b36416be9cf05aa5cdea3f977f46fa1c18a3e9c914853d2c2ce1ec84946deea32fb90975c2534ffd9df5312e8288f28c3c0a0a1df00091a65dacbd15e9328b0;
endpackage

package dat_33;
integer pat_num = 33;
reg [767:0] input_data  = 768'h680f66ce7176215e818073cb25947f4801e7f774a73a170eb7985e47459883f944a31ae6a1b52af0df7d2154c9ce9f3b729f271d9b0561623a152bcbc9845632311e8dfcad6d84ade97d5a353b54f23d8857f92c14b5f6a9aed49dc1ec7cd7da;
reg [511:0] golden_data = 512'h25b9c7dcb3e834d2bd138a4426f085442add46c4eaba26d27c7f872aca6cfe662654e3bc8e6bcdc38d86de6eea7ed37b85ca282a84021fa07962046dac1bcef0;
endpackage

package dat_34;
integer pat_num = 34;
reg [767:0] input_data  = 768'h56df7ef552df93ad321de58330d27d28cd36f470d1562161f40b72d5663040c95f4c8b7c51bffad381d819576c8a569419d52c83b8785b0cc1b670e5daf6ea965f20bcc0f9f82cd752370d51dfb46cec5d3161b35bdc4d4b5ea91ab1c7f7be20;
reg [511:0] golden_data = 512'h22e5329f4c2b9d7d2610fecb4f5b423b07b280cd812fbbfb29709b2bb5ebd37813ab6ae5773b8f6ebc05ea6fbf4b6128769d25261ac78066f896bdb03ae95e02;
endpackage

package dat_35;
integer pat_num = 35;
reg [767:0] input_data  = 768'h565dce43a31fe29b51a87dd3fa8b684bbb7c5c270f661aac54efc19b44b98a4b3b3a3e39e1c91657ef87e2030081dfb5f9a707bd3d75f5ab8d450cf924e8035c3ab6adbcf0b73a59c50d1d814ebb9e2c122b42311719bb08d02881cadee674be;
reg [511:0] golden_data = 512'h59f0ad6a684aa5b735537a2f45fdb76b0851deffae56251bb0ed669030d737c65b5402fb84e594b7c8254983e4f3e1e42b44f512b06f2b27637e4335e4317d20;
endpackage

package dat_36;
integer pat_num = 36;
reg [767:0] input_data  = 768'h5f781fc7e02f6fe737fccb5a494f5ecba2a5b2ffe59de295a3b278012da6602554b1f00159f0614bf37e7500998e7e02946aa970dba2cf5d262556458d3a6aea26138deb15a36fa84763a97b48b87b5531087c9b1d1bde370ffe69e528fc79f0;
reg [511:0] golden_data = 512'h19968ce551692a9c2a475069fdcb5516df2a7fa2182e6964f4436b7892c1779c4ba775371d00075d2afa8dc90fad14ee245066f3d270dff89459a91e35d73f98;
endpackage

package dat_37;
integer pat_num = 37;
reg [767:0] input_data  = 768'h3b61f91436736bc3c092484271b8a0cd587b1af7d0c553f86da9406f39abbb252928f9861f6a5d7d899ead31d1b09fc8320acba2c526361d32f38ec00d737e16476e1997e29c577a38bcbb07e9f42808123ab8a4c093d8796bc59d1c2920b70e;
reg [511:0] golden_data = 512'h3ee2cdb5fb736ddab5d4eba8067be937daaade228a5a4088870093eae5d28a54499f52cce24e86fe3043b4d8be96a031c1f3e33e1c8a22d732c0d5668fd0ce02;
endpackage

package dat_38;
integer pat_num = 38;
reg [767:0] input_data  = 768'h61c10c4c0c7406421ce7e91c738ad2c9a939191ecbc1a7f949a7545c63bb65e558e1181e4dbce4fd37369380f920777cc32fa2bb8d059bed0dd33dfd3e1ed54e5032bc95c343d9cb1af918d03000a6443e077f06c74c952e3aa1ce336bd0fe0e;
reg [511:0] golden_data = 512'h2fd02bcca8409ee391596e0669398324cd1436829c6bd9942b060813537ac3fe4c2520acba69a2af6c13d7ade12a7bb8a4e50f5214bce00ba4cd47e770969002;
endpackage

package dat_39;
integer pat_num = 39;
reg [767:0] input_data  = 768'h499bafe98f77eb7327c5f933a44cbe8e882fb6b6f5b87db1f644456a58d5ddc13a06647b4f8d8b6d171fc404441ebbff067df8bdcd6550b80ab27cf58f429e3c7614b28056d50d4f38a07e7b344402b58e34af558f2c38328c7ed41a42aa6fb2;
reg [511:0] golden_data = 512'h1c44b57a3e94a8887e5aad8c6de3a4a650c7fbb3a124d2589c1dbfe11c92a9b67c9e8adc6e5cbc89fabed909aa57e5b0a17868f12d5a20bf36de028399f0cd92;
endpackage

package dat_40;
integer pat_num = 40;
reg [767:0] input_data  = 768'h2dc0c7b1710ad550737581250487e0fe3e0edabf5551a94ab090d831cc2448d77eae80cc9e0011d2dcd74a62787695581d13de9675f60d43adff2ea8b5b4eb5e53b53380596d718c24faa3b680d222548114769fac1611e543f75d28de5d3552;
reg [511:0] golden_data = 512'h45d74b9f5a8e89c52b4de834f88f5077b2889f3f79f63320598c8953c24e386e01605ba1f0f34a8ea11feedc2f70f2f206641c2a511ca9ee56e5596f9944201a;
endpackage

package dat_41;
integer pat_num = 41;
reg [767:0] input_data  = 768'h4f540abdd5dd9fa8fd42dec02dfe1e859f03732a6d2d7f574b5d38031dd364e81d461229ba63fa4b6225c89808bd3c0680a9d83c5b5fa336ea1ddcd1abe282ca38d0e8e13e0b8a591385b887806b49710bdc4928eb6aa8c337f431e2f4fb9f5a;
reg [511:0] golden_data = 512'h33c71aab49f184f985dfbea85eaed13c5aa0114e872d1494115e1916181006d8295d886ffef9b0719d8770f87a00ac42a7da3f71743789aef6297c6584c4c2f2;
endpackage

package dat_42;
integer pat_num = 42;
reg [767:0] input_data  = 768'h642feb66460ca9620604e8f0cefa4afe000e4ed0bcbaaaab1c5f16c02dbc6a9432ca2acce99d8f388ee492f1a2e0c7c248e959fc59411bfa401feefcde45d904169207f5d9424ba6f246f17a04c7957f162d0cffe70ab433ca65732de33ce696;
reg [511:0] golden_data = 512'h712d78cc0a828447a1b3df75861d6add320360a9b6df5a0a0dbc6adddf2cb1541f104d665558f4695a6e0fc101ecda1653fed39cfb2000d0520823d6b181f604;
endpackage

package dat_43;
integer pat_num = 43;
reg [767:0] input_data  = 768'h5971fc9c1600a746d38c79125f0f7acb24ea9d7afed7c8034cf81714926b5c7f303c76274dad6b86cf5ad6f098d396a62cf75638a899d83e0e0a7003d31c5e7c2e8ad3b5cbb0c250b1d2c68942786d063200eabec3b647b4e76c5f68b9666502;
reg [511:0] golden_data = 512'h1b8d6428af57208f2ffebe2692e13aa029e34572343e9a93ad3d4d17bc43bcc268542cf86c92719667587e21f531f26438ba8f4b8aa6680385894b349d70be48;
endpackage

package dat_44;
integer pat_num = 44;
reg [767:0] input_data  = 768'h296e8c393ed3ff060645d5f398be3d43c55d00b4c57a615dea5818c9045f05c75b2218e0d69bf4dd8c6c7b00bd780184ef563b3048e7163c0fd1787606993e5e7ba5b7398770078b4718cd106665635071deb6f7cdcd9f2c1e1a30578023f5ae;
reg [511:0] golden_data = 512'h5c47773ecffa6dd5d75fb23724a01dab7d1925994fd9238871d9da64d94c80920deb330807deea243fbbdb3b6cc271ae42c6b0b7f5b77aecc7419a8ee4f9499e;
endpackage

package dat_45;
integer pat_num = 45;
reg [767:0] input_data  = 768'h336c944974d2ff377a84f7b5dcd6ba85cfa19dd49a74f4205f2c62efd7de4bf945d25ae3886a335f1c9a3fb0a5952ba8990c06884c457a305584a33f107666fc7e0983045880c7ae6130dd23cd112339164ebfd1a03aa7eccf37242882a0308e;
reg [511:0] golden_data = 512'h3f076486cb61197a4ddee836d3a320b96e83f971622be4363caf3dc937b2c58c769594f54dca1d8fe956a7c65d4c58fbb22f237300a507843e08bc27db65b708;
endpackage

package dat_46;
integer pat_num = 46;
reg [767:0] input_data  = 768'h481db717b37391930f581458c5140a18b82cc25a694f2fb57de6fac9c4abe38066e5f6e2711e47be961fe13b30a2ee2d146ee0e2130c0afa14f836b2dabbb12e0f72f7060576ececbca6d94ed9adf35969e7635f2dee8419ef6be363d3c18a86;
reg [511:0] golden_data = 512'h74e3b62591fa571e8d7baff29f7c1cc612f92af766ec2d92185cb12b8c85c2ac46c2bf50e56780460f96cfaa9ace5ccd552ab51a104603fd4d0f6f1768c8342a;
endpackage

package dat_47;
integer pat_num = 47;
reg [767:0] input_data  = 768'h7bf4b24d4fadbed007264e1042979092245d1b43d15f2d80b7bfd16f7619cf4f7a86acf44bfa27c3ae07f94dae513ddf34068fa0f9910999808f98cff28cf8027705a290a5864b13c6247449c6fc31d94bd84d9ccc2a275ae39d1310678b5fdc;
reg [511:0] golden_data = 512'h1ac83a9647381fa9dafc3951d43f256d33255b571892aabad9a3649a23fbd49a5dcf41127912a5939ba0d7182232c1943abd1028641352b18f4c3f5600b66158;
endpackage

package dat_48;
integer pat_num = 48;
reg [767:0] input_data  = 768'h77d40898dd9519a2f904a346330c7f0de6ba1a7f3749a46910bf8937ffa14ce8626acc260020256c695be91f8c08117391028bd9c444ab0f6ce8529439e618c40872a885217bddbd99d724a5d64637064257cc7e2a8e0cca8919353653df4cf6;
reg [511:0] golden_data = 512'h5f547b9412577416e550de9f72b2a681d0ffa56079de3b37bbefdfd58c44480c4731e81df4b8baec54b85423c96fe04d1805a5d9c92e9c77e329db43356fc24e;
endpackage

package dat_49;
integer pat_num = 49;
reg [767:0] input_data  = 768'h4054794c55aa68471773625098451d860c9ea43ba6ee3abba32075b5e0f02ed5056646438a96c1813ff046c82c5e6c939ef74d56c5bc89d1098a7a99b2ce15e424852a13e6ee7ff59f9e46a3091cd5c4d483c8c12006e26c2ff5a8116a7519be;
reg [511:0] golden_data = 512'h07470bbd387b677bbc5c5e32e0d50c5230add5736022bb0721d6ebc9b8374b42156ef9433f5bf957a1a8ec574a34c9757bd8f259aa2918554cffdf03b23403b0;
endpackage

package dat_50;
integer pat_num = 50;
reg [767:0] input_data  = 768'h3e4f9c060da444eb5233b3c0d2b83b1581e70a668ee22eb84445f7085a4b925726341791793a8d0a60bbd5805df8acb3d81317351f406623985fedf17b4106562dd53562e311540c329a0d8eeeb779c7b675aea511a0b203b6cd78bbe3b24694;
reg [511:0] golden_data = 512'h005e5c2d354fbcfdb0c11451ff2fa694d72b6781d21e2b8421add0ed128138a662aff585efb556decaa7b2e23f60809f4d38d9b96d650d5d8d5a85a192bfe4ba;
endpackage

package dat_51;
integer pat_num = 51;
reg [767:0] input_data  = 768'h391ad709c87f295adfb351ce346a54d33a8a1f38bb21a8cbdf4b1f73ec3d80ef545c6cc4d9aa64be5580a56fdc6e07c5c4ef8d6b9cc9af0b539fd61d8c1ae5fa0da135afa260344fd07194e337c6cf5305a24734afa335705898748f0f7b4d52;
reg [511:0] golden_data = 512'h757b5f4a74defcb05dd742e291a90f194ce0cca47cece2f63789516d47052ece31b2fc16f97b39048df11d28962913adfaa628d0717246688d9f260f21f3c446;
endpackage

package dat_52;
integer pat_num = 52;
reg [767:0] input_data  = 768'h242df5abc33468d04bf963d766e6040aeea80ce24b16a55a3cf47b0ec19d82d902469760ee59e70f58eab3513a96b4d8e82efb3659c05e10961da3c61027b7462ed2cb013d247991486c2d40ae9b0b19675cc8521220a7c99a58f3c9e2842c1a;
reg [511:0] golden_data = 512'h09d7aeb0f0b002ea01e4ca36145084a673dbd1386324a433e526b042ef5a964419518058403442592efff784f1ad0b9baf044fa1765ebc52361c480d36dbf10a;
endpackage

package dat_53;
integer pat_num = 53;
reg [767:0] input_data  = 768'h5d63709af1dc1dcc8a5d285aa8fa6b11586f98e340245002a2dadfbb5e18b2ba7eef87a7895c8cd87706057d0befc7954ecc31d938a3654548f3a51ca16f1a200c9401ce4d354e2df4f969211097a83cc9bd201a8d917279c9acd92b4e936172;
reg [511:0] golden_data = 512'h013de9f2e045ca40b1b5fb1eddbf634997c50290cc9f522047a756b8cbd23fe260701e92bdd5676f84f117e26b75e163ca1d0277b7977dcf9fb49b6aaeecdaa2;
endpackage

package dat_54;
integer pat_num = 54;
reg [767:0] input_data  = 768'h553c3709fceb67bf5896a2f382697dba295a2df6f9cfbc3f38c4020ea04bf15103b7de9ee8660f979f66846a3f9700f70f32aaeb4e25da03f9aea43589f761c21766e7f7614e635829ace87e2d3159445fb51dd14ad2ba26844fbf7ec8db3ad4;
reg [511:0] golden_data = 512'h7e3f0200a0b9d3bd9745fc422a92dd7e7c6f5608af13c58ea2fc5a5ad8c7535806e81b865fbea39c5e9f11240b75bf8cd3ef958134d7d1b5b8544a75847d281a;
endpackage

package dat_55;
integer pat_num = 55;
reg [767:0] input_data  = 768'h34293e71bd3b237b0a0624d72b597309f6d2b2d535cceeb9cf34a8e5a746a2f5225e4d05635981ba3b7a55835ce638a138d02c5c154168d6aba44f9349cd6f9c500d5af3e78c1b06fe883944edfad8938d994d0e82d49cfd14fee8c138f52062;
reg [511:0] golden_data = 512'h3f71d2f38428ea9d976607cde92949b4fbb3be4b28ca6b33ec6ac9dbae5f86584e1c005011f732d4f552d5a9be296b95908999eedf9dccc8928b8db914e9b5e0;
endpackage

package dat_56;
integer pat_num = 56;
reg [767:0] input_data  = 768'h4aaae6a832ccbed7703b16c8e9fdb7e31cba2bbdb28e53402ad97359f2d05581182572a3410a2eda136c9b3cbbadee2b98d627b0be29276fc7bb898c297998d863ba98ae4f8e215c6af34b85e243343acf9d91135d555b3636375ea5aa0514d2;
reg [511:0] golden_data = 512'h521184067ee448df6a0f74e415dfdc8fa4cf9d352624f9616ebf1524614821aa6ea136afac44fd679bb8075409d98d228aa40522fccb35cc4882bc178b11acd2;
endpackage

package dat_57;
integer pat_num = 57;
reg [767:0] input_data  = 768'h6b2a06eaef36f5ddc00da4c4ed61b3ffe3132ff65c402948c2ba6aa48bded1ea23932b2ff218e5855b22cfb7f89b0a02c3378189c824c3a3dcaa60dc6bba695263060a9c944b7d5faa08fdc48bdc3ce0a93b42d2a37a6d120b973bf250b2b132;
reg [511:0] golden_data = 512'h178bba5653a9ff82e88153415934b1f337f93b0ff59212de3e27d8c353b9dd760f12bbd5e7412491a989898dbc7342cde5ef5732f8af980cf59803086a134714;
endpackage

package dat_58;
integer pat_num = 58;
reg [767:0] input_data  = 768'h51229b2debe6596f6b24a2af4f608270c0f2234727617f210647d824f6eba9433d57da61c6502f5ebab384bc233c68c4d9dbc104c8aded8810080264d86da5326256a25c9360f5f6a2860082e39db7c0b09e13d94ce43748ba195b67408523c2;
reg [511:0] golden_data = 512'h4f22456994dd1dcfd87a6e699326cf56bab21f5bb789cc444ed5657dca6aaf0c7568269373910af2f992236789b461eed3861065b91232cdf25ed6ae338ba2d0;
endpackage

package dat_59;
integer pat_num = 59;
reg [767:0] input_data  = 768'h2c352b2d58956e6db68557ce3e02e282f364f7c989c629be71fdfe3c0ad2b14a313101132737bf31b77f6d006bef9d3be34c26a44d6b865ee097f0951affabf202bc0b8b7de568049461959e476ff0197804740dee39bf456e7eb5c458bf9996;
reg [511:0] golden_data = 512'h610374316f19b34800f543e200f7318e8f75ed7d5e7dc4d7e571c302bd06ef9c19aefc20bb6679f2601c1283f410f0de3347a763e46d5d20d01c67d9765f218a;
endpackage

package dat_60;
integer pat_num = 60;
reg [767:0] input_data  = 768'h01d78227e81242b848e10b1846f3d892ff8a656cab7d16c34be961ce28e51c20247f7cdbd11a0bde55855a463a2201a1d945253ab36d10b38f871049e003a474350736526d0b725416291ad2699f4acfa5d3794cd01292d4e34b52acded92302;
reg [511:0] golden_data = 512'h26366ef84237ec542f18cfd2b7d3ef0bb3ed34b003c92448ad292a12ea60d4ba2eb3e33e3f41279af0b93215514708961208580d39dfa08cb78a323173485052;
endpackage

package dat_61;
integer pat_num = 61;
reg [767:0] input_data  = 768'h6684ac8fd47b667931f99f017c855b187db97e7c817e2bbcce8b1d96fd6f26545662d31c10684e3ba9f0d8e43ca8b8dd50d6c91d563c2e1666e834172dd5f9fe1ce7687c2f0d65fb74d73be223291dc61916967ae9f736695d3b9d39595594de;
reg [511:0] golden_data = 512'h0b4d1a2144081e20a2c2eab7a3b7bffe7c45a6a09cf74d54127860e5887da228735d77c5bd853ce291927337ad29785e6e2321baa435631effdf7deff5ae9944;
endpackage

package dat_62;
integer pat_num = 62;
reg [767:0] input_data  = 768'h4fb24b7bbc78574883da8cec5a753040996b05e570e0764c461cf72bf516d33e5bac2cf683bc3a8716b50a6bc299b916f051596dfd01994c9a53d287f5c2ea601629fad980fd8e592d6374a7fca5d7296353357958a1ac96d05a9e5d038673da;
reg [511:0] golden_data = 512'h0023a396ada1d511581507a6f3c42314e90334732fd476fe31238cf1fe216e5c17136d6b91bf0e371092f09bc34d9aca0097ad9b12990a355d47496389de83ee;
endpackage

package dat_63;
integer pat_num = 63;
reg [767:0] input_data  = 768'h410b5fe4082f1be4d942ce9bbcec2d076775e0275b930201cbf4e547b0fc806a587dce40e6473052ea867e8fbe2d339b21fe6cb59163a71f045c945e5ae5add226a55968896daf409f6cf8a3b2151c0444d799b0f377320d8d04a2a0c32dfb54;
reg [511:0] golden_data = 512'h677b0ad2e1c34f20d51401c8f978e62edbee60a72ea6b1247c09fbed7a7c771e03bb06d4e9dd22ef98b15b14ec25eb663a9ca3c162a24c45aa2547d34f60ee7a;
endpackage

package dat_64;
integer pat_num = 64;
reg [767:0] input_data  = 768'h19a0593ac8e26c60654d387d4c7dfb2bb26855026c179fc9c40811a2e62fdde6025f258e5097f5193820961f9f0a6f9d0a2038dfa0d64a1e95b13fec92d3d1c020ecb31bcef9a7ce94fba5bf0bd8150a56770d2989a3c2db4f8149c8687184bc;
reg [511:0] golden_data = 512'h0231949c64ed9a3dc617d1e6aeb68f21f37c0dd0a43ce92e6e3ea4dcae1407b639dea66e86f7bde262aa8195c7ff08152538e6893031f1ee370ede0f27607056;
endpackage

package dat_65;
integer pat_num = 65;
reg [767:0] input_data  = 768'h5b166de544ba14c7e1479ad2982bccb08895fa92b1599ead9becd744bb46846d12e7f48e2196501ffbcd4876a181664864040af139e2e419e1f21c5846ba959047bcd965379b369fc0bfa7723efdb846a32467a1f319c28f894938c631718068;
reg [511:0] golden_data = 512'h634b92bcb51c2e6c52ffedd7f4714d19ffb9351c87ac901cb036775cff900b7279646fbb36580394e6046e115bc59c990179a9a3ff6e7079d58820589eed5e9c;
endpackage

package dat_66;
integer pat_num = 66;
reg [767:0] input_data  = 768'h44e5a1d3f6a7b3e9f8bf2547af45f148959e5eebc1ad0890e98b4be71e1fabe410d5594536f9322a163cd795f5cfd59c08c9fba176d7c3852cd949709445371a35bee164eda810812b606ae58cd740483b1bb699a0ac6fadbb6984ad548469a6;
reg [511:0] golden_data = 512'h37962a5b11d0be27bb1ecf2bcfbb2f27d92bfc78b862a850dfb296e6c1a08d4004acfed7ae4c587797a3c454791aa27251cc623e533cccd99923c2f1cfd07548;
endpackage

package dat_67;
integer pat_num = 67;
reg [767:0] input_data  = 768'h4a1c98d137329817e5b5dc54d170edc6a6e5cc78d2e98e4777322572fa9be9af4aff72182d7a83ea27794960491b9c20b06d5500149032c4bbaceeedb6ad7a985edd9e767675e59ef143e4d38687943e0b5f9371a0b9345ce8393c9d5340f98a;
reg [511:0] golden_data = 512'h4ded8ae7edf4b4469fa7b3d36a0fed0104e1ebd522cc8bc5bc72af34471f0c7e1ed31eca8bc2aa8a0d7b6ec300e1377771b6ef00dcc7c22154413358e6d68e8c;
endpackage

package dat_68;
integer pat_num = 68;
reg [767:0] input_data  = 768'h4ee9fe7a541cc454df05ace1c83eb8625a4296930d5cbf683f6efe727cd39e120fa6388dda177fa4b43397dbfadaacd87806e3b8f2808cfbaea4d66582ca0f7819d264430e4cc91adf82243ba3aaabec45a5610bf5a9373aec72fdfc034d9138;
reg [511:0] golden_data = 512'h1c2931157b75951a6709c4bc95a74d6e89d79629d6e685af9d06759c7a33c9aa040bf2da4d4fd3a86bfad740c9c036259aac2a9ef7a24138b644ad636ac5ef52;
endpackage

package dat_69;
integer pat_num = 69;
reg [767:0] input_data  = 768'h3991121df09bcbbc54ab64e76c5e5f643af27f5d1d5d6c3c4d86b88a65536d802bee4e68e62b17121d5f184d236c6b83fe1c92f97cf5bdc389c5e1018e7210d05c5d7fd5d4180b8bf0d47ef767c8404ca07f57e0ebb0e2cee48861c11d3f2568;
reg [511:0] golden_data = 512'h17a25e86e702c4032e57c008b67bc7aa078edfbe682cf3cbf6bfad55ffbd798c551d32f8cd563aef1bc12dfcc70297cdd9d296a57f01f03ff7dc8f79c7ecc94e;
endpackage

package dat_70;
integer pat_num = 70;
reg [767:0] input_data  = 768'h57f9058076ad04ff63751fbd4488b0f51ef794bd467f364b63ca2c38a7ea9b366c67dd9ed8feb6a200331b8380c8e0f77549f9dbdf346dfca1dab98b7fe3c654042d5032791b17f2fc498ea71ea60c809b59b58e3d9e2c722901ec3864daf07c;
reg [511:0] golden_data = 512'h16f73a7c1984493bde060b8ed4e513b46edcb9496e90f4a73b175288197d6c0677c153c06c09e3ea1452892b87d1cd59649f25df89a991af33155483dbde4f20;
endpackage

package dat_71;
integer pat_num = 71;
reg [767:0] input_data  = 768'h71ec06400ce34f4f8f9635a6dc9fc56b71e1d6d2d44fd0a43471df27a20ce2267e5bf703991fb190426ece64f82fa71c5893f38a13b225cbf5fb13dfc5db3a7c276b23421bcbe96b9b9be07f543f0827200c32cef62aea78e23bfdab21cb1d00;
reg [511:0] golden_data = 512'h45e2c06053ba8f8916bbb82550178d9f095ec15bd8fd89f0f1142b0f2603d1f62ee12c2f8deee756728fb73792515791277572b763c609d7235484242c05c09e;
endpackage

package dat_72;
integer pat_num = 72;
reg [767:0] input_data  = 768'h08a7a7a50d92d70df003541f60c1f1d59574e76484ead36c52f1ef8e14f854860fe4f8f8cc31943f7433d651bcd947a11a262218a0c8650a5280dfe522368e247a53fa00ab439816ffd65dd7e34d2c1e1ba57bafa06630401c27b2c23fb6d318;
reg [511:0] golden_data = 512'h536419faa722214b07a5b125c8787d5d72a504deb6768ff39d44df7f08e060826c7a86a5b1336592063115a7ed657cabeedc602ad4e30fad1ca24793a4cdddaa;
endpackage

package dat_73;
integer pat_num = 73;
reg [767:0] input_data  = 768'h47e79e4e14164195ab1eefa72309ab5d9e55ba08018b7a40ec287bcec0fc00f37ce362e4b61ea8c7a661b1ed70f8205ccc0e4ef880bd30c57002521fc433d2fa75384000c741d4dad5371265eb86016d59f6e446db9e13e2e5252c90b8a0d0c6;
reg [511:0] golden_data = 512'h43e12b0b9dfc7a199e38e17a9465ebbf808fb01182fe462b59343ff040df849e3827d1cab85bc09eef2497bcd91df9542920ed1377d0fc1611f76d1151fb9fe4;
endpackage

package dat_74;
integer pat_num = 74;
reg [767:0] input_data  = 768'h7fe2c687041b4264e5490c39356b68d50d6fcb2adacca0c4324afe4bb4463a9431d15d0f491f7ebac0f343979721ddc181847133a8a074a4443e634bd3b2865279d0a7cbda89df89ff1639cec1e067e6caf9c5bb6184a6a4537d35f0393ffb2e;
reg [511:0] golden_data = 512'h22060aac2604275786c5039a853624d99f7033cd1581ef2083134e1083aa98f23d9af35495afb1c144fc7b661188a8d179f7197ceadd921c378030f732f7eabc;
endpackage

package dat_75;
integer pat_num = 75;
reg [767:0] input_data  = 768'h4211a57b74e57f900e950482d1a6295aee10ca705769086f5fd3e814f526a9e16fb4f4793f87d3fee658b256a5347680e516486648b39f30b00f7f7cc0b3395a700f9df2053d07a105a0e858cf6f070b953c97ca5b1930d1b80df3c483c1cbcc;
reg [511:0] golden_data = 512'h2f19ae95c8fd45180619a7df9f3647c34a7ed02a55287aa71c004ce9a98f04ba37c7653937f4484d48db444f8b0bb6ea2fb33b0d3abe0c2eec95aa61ce378204;
endpackage

package dat_76;
integer pat_num = 76;
reg [767:0] input_data  = 768'h59f04538c9602fe125140273011e82d124687ba56bc1a20dea75f1a8640fb354119cba15bd93e5fa3168f911dd65d953ed9c9e8e28aa3c827e0824e51b06b1c667ef9348a89fe55b6ef54344eb303bc47c19f3f88b574c8d47cbd20723dc9866;
reg [511:0] golden_data = 512'h2710f57a7b16047d6da3869d42d90bb7816ee5a251287669c88af0357a6372561e828da8d06887e18e0abbbde82210b0afe04ad5e8e1401876859dccc2bbac64;
endpackage

package dat_77;
integer pat_num = 77;
reg [767:0] input_data  = 768'h7fd88826323f166e8148b519ba62ed3a0771b7f741cdf885062fa234059e945f7aa558256c77d25b2e2916e0176bb6cd9ac0c11b7f32ea282a6bab4ddd008380254f84118324ca39cb04d87a0c450951c54539ee201d638d56349cbda82856da;
reg [511:0] golden_data = 512'h5412d335d34d30338958e06266a8f5b3a6761df0e49b4d870cb1479c859110a830b8f1857eae3e5822933e5aecf9b81e953167893aebc1432daad57002c8e0d2;
endpackage

package dat_78;
integer pat_num = 78;
reg [767:0] input_data  = 768'h71e71c3cb0cf01a80066002642b43160166bddf43a92c93b0ce58781510fdd0f3a471c32d0fc54c85eeee64107512010800792e7d9490721c230f490fc32b67654cdb7f06e0570f47c6c4a762aaeb68da98abda2cdb133cf6565317a39c29216;
reg [511:0] golden_data = 512'h72aaaee6a0d1c0024ccf7a408e71627f7f1cecb9c8bf406a42e0e6336cbb7918020c2c5f15ce87e6c3de58ccc85c4261a7d5d838cdafd5233cac2c584ac198c8;
endpackage

package dat_79;
integer pat_num = 79;
reg [767:0] input_data  = 768'h4907f18246299fb2141ee10d28ff6a5d3d70add8d4b99cc97f2c39ed970e7f9629d226dcf7e880488c9e87ab5a8dc698d551ab15a3c3e69c86cde53eec4f87c878cee2b9f7b9d44a0a3b0cca72d343ecb9f5876c0fc03ba127ee03e30a25deec;
reg [511:0] golden_data = 512'h2dd32d5c5eb80962f9c07a05e7589f77b58bac95179e8d965ba55619189e8598684e8386063cb1e57b7599e1ca23993c32dc5540bf642710340d4045ecd717a6;
endpackage

package dat_80;
integer pat_num = 80;
reg [767:0] input_data  = 768'h5b2515ad94102be4ae5251d6a60f8eee04ceb02b1fbbe81009115a34e58c5e5965579a3cac964fd20c495d179d87fe0ea1a1c18a9f474c32ae96845328abdaf240d4c7ff6d49d963bfcc724e736b40e4fba643877ce9a7a7207da5158bafd2c6;
reg [511:0] golden_data = 512'h276a0fae82673752d0d2ae48d8c316d99440771b38066f68c066898600a1eacc2c905963f5f42dfb91aa075fbd533a745b0a99360af5fa02af37fc6b444220da;
endpackage

package dat_81;
integer pat_num = 81;
reg [767:0] input_data  = 768'h1a0e28f1c400326e8dbbde9d3d2673877c6a4e09fd8daca4dbfd1829d0e803df232e2db035ea0d6cf40cb7c7d75e9545c6fd29fdaae5944473b307ee8280247a1e93d0ce8d0a9e7596eb303f12a39c79af55cae131340ea8c95658d95ac28fb6;
reg [511:0] golden_data = 512'h4180fc9d15f1fc23f4ca385511540023af2fce70561c51e640c05258b082c2b6289c5c902f55ebb9c36ab2be4997e494d6a9f13e9f4f97b4f419d24f49529602;
endpackage

package dat_82;
integer pat_num = 82;
reg [767:0] input_data  = 768'h22968de2b67bee4d04edbf06805a0b519155f24ccbc7628d388d5aa647026b3748e0b5679c49d45d7a78f9e58bfcfbc402bc00155f854f1599bd97b00d5e1e3a6608721a8c5443e370743154ce74f2bd780b1e9baec947a3b87e3b9a8e403590;
reg [511:0] golden_data = 512'h122739d5a5833a74018764a9051a62864cddd3e3969ff28ebde298acdca3e1983907162eacf4dde79b3c0b24e7983273346062587b758a4da8e740cb5aa1e0f0;
endpackage

package dat_83;
integer pat_num = 83;
reg [767:0] input_data  = 768'h73c4733c7e9404d9841e20082c34740bb46ecc40c74b846a6b9b6a9525a508c617cca15f1029ad93888d52a742144c1ef3811bc15f8582ed63edba1792febc1664f4776e8fb3526ab7047ea5bf1c87432ce5e5ffc66909052d4bebf176f6398c;
reg [511:0] golden_data = 512'h137bd57bc2e0b006f46f07a5e7068ebdb33148ffe36a7a9d1eab70fc83d7e16c7e64ad2a1b42576801930170ba9525a740c1722cd86c3d76abbbc8fbb2e70a72;
endpackage

package dat_84;
integer pat_num = 84;
reg [767:0] input_data  = 768'h60f35d1b91603a60fc39caacf5405e050891c2c32d1475db213b5e734b5a72db0f79bb480b968e517b07e96ee3fea7559851b7577b9344f864614836ccb67e0c3ce678cbc4b1be70ea44f1bf571ba1e79867cf9f0546b8a97a0274854024b1ac;
reg [511:0] golden_data = 512'h3dbe3707a0912859dc402df42eaafcd63f130377bd26ead6a912ec9e90a7fe4a699206b5dc878cf8587b39a70ac7f5becf2d36a784eb25e90e5c33da9cc29608;
endpackage

package dat_85;
integer pat_num = 85;
reg [767:0] input_data  = 768'h02e84ed19d33ce9eb1e393733c7e7a5377e6a4f21714227474d6b2f658cad33a613b58e30b62d1ee671a6c18ca33fe55992d510b8b6994d7f755f28d6a66b1c8262db067f8528f4ef50bf0604851a71cc2edf4c60f843fb3fe9fff27ff3747ba;
reg [511:0] golden_data = 512'h6ed0ff4604109e57545aa18b15693579aa9a37c6fad900bd5bf52027855c23f65417d02bf17319a97023d8a67146e494822f747e77b9b54b05e073a271f27636;
endpackage

package dat_86;
integer pat_num = 86;
reg [767:0] input_data  = 768'h229098565eb0e339279be511bce9ae96b91134c16e7630845f60cb8633a23e1c63fcd8f096e92b10710423322a6f962a5530caff0c830a226877a8670dc6df24614a5e14dc6bd37c7c7c9ff018d3aa3dd6ffb9cdecf4962db6a96474ccb3a846;
reg [511:0] golden_data = 512'h13242757572156ccd5a66abc773cd81d84b3d7bface9559b1af8fe61f14f767a3c55ca93536cbb8525eb69e1140c583f2d7920838998a65da6f4c9716093f634;
endpackage

package dat_87;
integer pat_num = 87;
reg [767:0] input_data  = 768'h543e8d66ae8bb4879699e0abc2d5b0598cab80426644b863d655114e2b3f532d6eb0b771c184a7803e95c30d7afc62520bf4863019e406e4d5239b474eeb2b346df34470fd6a3e9934860453f7b9e3e19f6124c0562c7e68c13a626c6d9b67f6;
reg [511:0] golden_data = 512'h46d5634b30b38e574b3229d9ce00e7efb20b2a625034febd9916a3feee3ad0ee7f934f11ea4d2719aef7fcd72134d742fa7d22adea54651b2ee0c95c74c1d294;
endpackage

package dat_88;
integer pat_num = 88;
reg [767:0] input_data  = 768'h74f285ae3af118f2cc70fd3e97e550524d07d04984c4eb1711fa0ac422dba65303a8d59573fb2b7025aa051afb42a8827dd6da0c0f454ae8a5dedb050f4ba85a4775235362369d6b73d4d3bfc71341e8394655b2c760e0511d53a642831cb4a6;
reg [511:0] golden_data = 512'h23f59112deecda02438d2471508ea2c7a0bda829a3cdb35cf8819ec49b269c540a7e1a598a23c821b572fc92cba459d96e863965b5db6ebc72b97d1b9e4de342;
endpackage

package dat_89;
integer pat_num = 89;
reg [767:0] input_data  = 768'h1bc97e09f23c0a9ec9d436fb1f91ee20935dd2d588d6ef936e116a6d3453b54f47c8ade9bdac925d056ae03804db7112e9c17889509bab1f8bae96950e30e2fe5d82b85de02524d13129fac05d51e7e28855033f2465458e0b0f426b003a93cc;
reg [511:0] golden_data = 512'h0dc9f1c842730a25db580abb046075c3c93b0a3632f57e1ded47b4b5af187b0a6d26d1342a89493c9f7cd9cbd23da6d46922c13b77f926ff09cff4374d8721e2;
endpackage

package dat_90;
integer pat_num = 90;
reg [767:0] input_data  = 768'h5c7dff78789a3fba533a6a42da56020ddad7749b44d40358e97be86b30b188871883b2c8cb9ec29e307f1c2ebb3008e25fbfa9c0c350f2c3bf405d11cf2902742312db8eeeffd3e0dd240e04037f6e6e14da91bb33ea9159366a30b27c9eef36;
reg [511:0] golden_data = 512'h5f6f5e214e892e7fc2bba217e790d4460b12225b8741299835360abc140b35f83e72379b7f8792d9eb3c227a7ac19991753594e2d7306008805af26c48b7763a;
endpackage

package dat_91;
integer pat_num = 91;
reg [767:0] input_data  = 768'h0d7af9d01857a741a571fa8bbc97d8bb5c787a0930b1e06754d9c75945c235d705dfae39be9ac551b25b0e9518765a972564f9e3741d9b55ddb56c00bdb23240635acb9655009086e1d96d4d57c7c2b7c9ac4a2ecc3a818937b8f578476626ae;
reg [511:0] golden_data = 512'h728a078b1652a9d9fbfee87345d1a5412f6612a6fbedc586c6aba4d78ba518124e98fabb575660f715d11fe81f1d5d3e6fb68d8c9e308d622c1221a621f4236c;
endpackage

package dat_92;
integer pat_num = 92;
reg [767:0] input_data  = 768'h4ad088c343c33d990e4d9432a1d510406eb6ddf0ed60103dba7e4c09305b195c0e6503241670a4c429660bd399ee11d4bc21e1e9b2d1e413ed7f75936369b9ca6b936af1f9254bb178f9eaa9c83bcad09a3511b8552b2917c7848f544c62a014;
reg [511:0] golden_data = 512'h48d5470ff163b1663e350ccd1e7195313a559e649113e8b97ff3eb6713e09e961a20ca1eb8f5cdaa4a7f3274fe54a7e6a08df44b775fe1a6cde99d91905868c4;
endpackage

package dat_93;
integer pat_num = 93;
reg [767:0] input_data  = 768'h4379d268c6b85cf40d353a662a64bb8a362046daf6e633d61b162dd57382bf9151e2acb1c50a2dee37db85ddcd9cba6cfd0042ae348184a50b5fe1634075ca7c3c65cec78f902be674543290d125939d83b5b55148cf5b474dec0e06e3154934;
reg [511:0] golden_data = 512'h6581afa7a4a9c4153d982725d8a82003629ce27585ef0fe0d45a29f9185e4d8623357b03912e1e30fb65f32b6b168d51d09e6b1dfc5cc3f791f76690337a44a0;
endpackage

package dat_94;
integer pat_num = 94;
reg [767:0] input_data  = 768'h45cce553c4efe389459f8ebdc2a939f84cd4e5dc6404f52e3a0338e0e004179032653efe6f02cf381121260a1903c1a48296dc54a04ceb01e94b567db7b62c406cd92f971bfd5d4b885e7cc4359e5906efef065dc14e1df2e9775483ce5d3a82;
reg [511:0] golden_data = 512'h4c9cb456fe86ff845e3d13217bebd11dd1ac130dc79c3f72950b2e9ae7d17786794949faff884a404cf3e64d4724aa71033e88c6f293e914497cd8ced0ddb512;
endpackage

package dat_95;
integer pat_num = 95;
reg [767:0] input_data  = 768'h378a48b973172b420969d1432ee61061a5b51ccebb6cef0463dcb97905ef2df77c9f35e762d974bdab6f141bbf90165b955b6b7f2d3e90a3a5cbae354408d7c61076d89ae77b0e2c9e965d12268a2ebee42ea68cefed3f7ea72fd8c62f3d8266;
reg [511:0] golden_data = 512'h58027dbeb5008c033949be5f5b6b99175a29c4faaba27da0283016a29c53776828430bb554facfe93afd089cc6c3bc15fc5573b634519fdad4b16a1e79365040;
endpackage

package dat_96;
integer pat_num = 96;
reg [767:0] input_data  = 768'h0d51cd41e30e7306daf287c9f531c1da6737b796ec713745d316639763796eda5b96ac844b7e59f7c61c1f66bd78bc49a30732b56e6ac640bd71d18c76a9ab3659b5e7cdba9ebe3c8f26c5abd8416f1c7b46eb0f1ec758ec52de35b379602670;
reg [511:0] golden_data = 512'h6a238a35e560399d148f0737f0b0ff223b42538cd37c5bb6ce7813106203c868352ed536d18f30dae2dbe6dde17415e07833cc21465b1f3e95518d84fa639f92;
endpackage

package dat_97;
integer pat_num = 97;
reg [767:0] input_data  = 768'h13606a5544c28b8b0e970057316a9a134e8f03025a21372a1580ae83b23b37737fd6feeea9bfc723878d82e092cacc838ae50c00358c1f1bf497aafc7948c102430c88900c64402e195c10f0f86c5b67a94fe6b610b2567a611de9f0c01ff046;
reg [511:0] golden_data = 512'h18c3cb496945a0cfc19de0a404f5e3ef87b9ab2efed3fa49a3bdb21b92cf0bca40a01b2e66ff20b37e6914ca0d09f23ed9b242f6158c86393d5fb61305dc0410;
endpackage

package dat_98;
integer pat_num = 98;
reg [767:0] input_data  = 768'h7cdd6279538457934f0bb63acf2a8735c765967cfb78359d1bafb95d504586fc0eeb86a89a251a6f943ae99ddae571f44403dd6d403b7e58c98a7e9f856d49347a29a75a41644cb9bef32634c0a1fc9046c66a3019cb54e679662ffeeb54aa44;
reg [511:0] golden_data = 512'h4c7ab3da61a6ac4c730a5110b244e4cbea22a3a3bdadfc3d58765b9d7e539d541726acd5550b99adca2878a77b99867486cbd75bf882e151424d5087e714f10c;
endpackage

package dat_99;
integer pat_num = 99;
reg [767:0] input_data  = 768'h6cb69a7975710370abf1e793c30cae6dbfcf5d7c593145229e2820067a1b10f07b8d291dec8a0c09a8b701070b7fdce9db338797c430ec0da06bc8f7c50552f00a116b57f9a00fa1bbd4d9809dd13323ce90dde78b9c51fe0c0fec6875ec0838;
reg [511:0] golden_data = 512'h0132692ecf282744e34587fbad888eb54683b9703b95976f3e9c88bd26c0c98a0d4bb87b8b52b1fca45ef4ee524d0219aacffd32ffb4594d6641245fa5167308;
endpackage

package dat_100;
integer pat_num = 100;
reg [767:0] input_data  = 768'h0200ce35af8709343ce4b321d953e87793d698c6e440908bf3e3211c128a8ab660131cc634eb4610368652b739aca5bfb2b184a481f214a9d390edbe5804932e1f0536af937118b4a58fbbf76f10ee19b48c63c7f8278354478f0ef72b4b0e26;
reg [511:0] golden_data = 512'h7a39b8c22b191eb3d3318b510125320b5e57dd278972eec52d55d54b43aaa78a2084a1e1d802685aeba66881fd0d866ceda2d66a2e3e5b1696f695fc76b5f0ec;
endpackage

package dat_101;
integer pat_num = 101;
reg [767:0] input_data  = 768'h2c2b71052d16b8d66e9a5f7a995b9b0243851dd367e6bb54b40977c5f03996ae49dd3c8e0dcbda66c1a632937a15385cb3d315733dc010e04123d0055a5f08542c38f78b72f1fc1749db4e2991921b5ba376ac8c567206cce588a64d438d8a2e;
reg [511:0] golden_data = 512'h74d8416fe7c5a2046c711b619a45a5ecd5ac845962578c116eb02d52ca0d67943f7e12a02662f3d220f231d38f47ed5f60fb8bf3508b004771b8050cbccbffbc;
endpackage

package dat_102;
integer pat_num = 102;
reg [767:0] input_data  = 768'h43a5b20387c3941935a6f273e0f105155d09bb131099426e7acb332059c9a4aa241ad4c41188b9ba2b158cedd82952947e9b636c6c18d267a03d73a76dd3d8622aa8c57a63c28ad3ed225500b135b2d2908522ade448f9d28688737bc79ecd32;
reg [511:0] golden_data = 512'h6f5e8bb4dd7e44d4bae15e28691a8fd85afcc2b75f019dfff2849f8b32c5552a639b76584650a84af3a5156733996a2b05c0f41181ad2e188fa6758cbcf0ebf6;
endpackage

package dat_103;
integer pat_num = 103;
// M: all0, X: all0, Y: all0
reg [767:0] input_data  = 768'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_104;
integer pat_num = 104;
// M: all0, X: all0, Y: all1
reg [767:0] input_data  = 768'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_105;
integer pat_num = 105;
// M: all0, X: all0, Y: rand
reg [767:0] input_data  = 768'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001cb76317ed6b7e5053aeec6a34289c51439af5241c10162118e7bf8ce3fa5276;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_106;
integer pat_num = 106;
// M: all0, X: all1, Y: all0
reg [767:0] input_data  = 768'h0000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_107;
integer pat_num = 107;
// M: all0, X: all1, Y: all1
reg [767:0] input_data  = 768'h0000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_108;
integer pat_num = 108;
// M: all0, X: all1, Y: rand
reg [767:0] input_data  = 768'h0000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6f946993d4cfcbaf423470ff3b32bd2d36e9b1d2c465541c7b51e1e80adbbd71;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_109;
integer pat_num = 109;
// M: all0, X: rand, Y: all0
reg [767:0] input_data  = 768'h0000000000000000000000000000000000000000000000000000000000000000ff4df5bc8a3c4b34be4ab2853e8c9e8420ac0c07dd28e8e98b5cbda2c94a084c0000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_110;
integer pat_num = 110;
// M: all0, X: rand, Y: all1
reg [767:0] input_data  = 768'h00000000000000000000000000000000000000000000000000000000000000006138a6360627178bcc404bdc5d5e9851c155012d111a3e044388dcfa037f3bf0ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_111;
integer pat_num = 111;
// M: all0, X: rand, Y: rand
reg [767:0] input_data  = 768'h00000000000000000000000000000000000000000000000000000000000000007f25cf27a452ecc097dd8afded29394f5f17b3ae650d19da0aab4cc9d9af64bc5414167f1bb38b6f63ade1e9b8d4f6fc7ac3f9ad9920f56ae4897c9303cde243;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_112;
integer pat_num = 112;
// M: all1, X: all0, Y: all0
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_113;
integer pat_num = 113;
// M: all1, X: all0, Y: all1
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_114;
integer pat_num = 114;
// M: all1, X: all0, Y: rand
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000000000000000000a1c7584939ae48375cc63ec2a84c036dbc5d286189e865754131c63a7859f08;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_115;
integer pat_num = 115;
// M: all1, X: all1, Y: all0
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_116;
integer pat_num = 116;
// M: all1, X: all1, Y: all1
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_117;
integer pat_num = 117;
// M: all1, X: all1, Y: rand
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0e8f12a2ec577976edafdb5a9c804813ae003dd13f1dd16447f3e46d2b2602b1;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_118;
integer pat_num = 118;
// M: all1, X: rand, Y: all0
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5f519e628ea004d5b09b44d627e5f9f9f5ba4c97e069432c3f87159298b81fdf0000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_119;
integer pat_num = 119;
// M: all1, X: rand, Y: all1
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed3ab062ed3cedef803580cb5212326d233829b4add68cfbe9a0015bca4ac98dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_120;
integer pat_num = 120;
// M: all1, X: rand, Y: rand
reg [767:0] input_data  = 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff508b351f2fffdbddebf670dea4f1e3e50aa5dd78d5540a51887d464fd7c7d97a8cf248f471143af21780fa063a4f581e2d80dcd9a52c02ddd82987abc46b6942;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_121;
integer pat_num = 121;
// M: rand, X: all0, Y: all0
reg [767:0] input_data  = 768'h2b0fb9f72198acd2a7173994cbc66b0770529b45f78f251857219d0ad28a7b2100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_122;
integer pat_num = 122;
// M: rand, X: all0, Y: all1
reg [767:0] input_data  = 768'h65cd5a2e05ba0bae9e45061290e76c08a023dffabf22c95257db2d014464c4220000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_123;
integer pat_num = 123;
// M: rand, X: all0, Y: rand
reg [767:0] input_data  = 768'hfc58264d76e87708527432ab126833aaaf3bd32bb7f0762e23d41b7e2cab6e050000000000000000000000000000000000000000000000000000000000000000472ec6c9422ea76564e6089b9cd1df92571b7a586f6cf300c183e59452f67f5e;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_124;
integer pat_num = 124;
// M: rand, X: all1, Y: all0
reg [767:0] input_data  = 768'h3bf66cba49e8dfc07985d60e1c3de91179b8ad8e64919cb2c78db974638b819fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_125;
integer pat_num = 125;
// M: rand, X: all1, Y: all1
reg [767:0] input_data  = 768'h2938a6e222a255afb259c93fbe0643103c2d76acd1e8a87c78e22357594deb4bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_126;
integer pat_num = 126;
// M: rand, X: all1, Y: rand
reg [767:0] input_data  = 768'hf5117063df99c04a20de9efaa2836273642238d2f5d06ea3430a529a43fde58effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0995c71cc56e9123b0d11f8ffb46c91adf8331ea1e9796802c184eb8e6a8a92b;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_127;
integer pat_num = 127;
// M: rand, X: rand, Y: all0
reg [767:0] input_data  = 768'hbcea55b3c34b3f5a64ed40b0fbf541ee822a6fd852bd86c85b3fab840517fab1b3d5110eba4dbb127cd57120854bdf8624d1c3110d3f6dbbe30a5c760d2b74220000000000000000000000000000000000000000000000000000000000000000;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_128;
integer pat_num = 128;
// M: rand, X: rand, Y: all1
reg [767:0] input_data  = 768'h7da29e9628f0dec3fe3a7908ac05ad2e702b5b578cad51394c7ca824d05ac6002015cf46c634940a0f5c3bc0b2e013104c529624d1f5ed8ac972abca9f7a302dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage

package dat_129;
integer pat_num = 129;
// M: rand, X: rand, Y: rand
reg [767:0] input_data  = 768'h48a6c1fe69b81e5fba16d584ae50f654a3a5612c33f392ab708752488b8beb3cb19cacfd123d88c0f716df7335630d94834745e4005c49ef377183a4567056abf7e9a0f83227a52c50fbc7860a2b26b36b24d99107b78cce2ae528740b44b0ad;
reg [511:0] golden_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endpackage