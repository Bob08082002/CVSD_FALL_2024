// list all paths to your design files
`include "../01_RTL/IOTDF.v"
`include "../01_RTL/Sub_Key.v"
`include "../01_RTL/F_Function.v"
`include "../01_RTL/CRC_Gen.v"